
module conv_windower_test;

   wire [1023:0][1023:0] airplane4_conv1 = { 1024'h003c002200000000ffdc0000001e0039ffed005fffde001000020070ffccffec000bff59ffed0006003800000021ffee0000ffdd00700032ffc7ffa3fffaff9100200084ffe700340023fff0ffc400190000ffcf004a000e0037006fffc7ffdf00000000fff70029ffb3ff92000000000011002b000000250047004c00140000, 1024'h003d003400000000ffb6000000240011ffdb000300390018ffb60006fff7ffd8ffe4ff8cffa1000900030000ffe8ffe00000ffdc00060037ffd9ffa1000affe80026002dffeb004700240027ffe600160000ffbd00820033004a0060ffc6000600000000fff40008ffd7ffe9000000000011002700000012005c006000190000, 1024'h003f003500000000ffb4000000260011ffd90003003c001affb40005fff6ffd7ffe6ff8aff9f000600030000ffeaffde0000ffdb00050039ffd9ff9e000cffe60028002effea004b00260028ffe400180000ffbb00850036004a0062ffc4000500000000fff40009ffd8ffea000000000011002700000014005f0061001a0000, 1024'h003f003700000000ffb4000000290010ffda0001003b0018ffb10004fff5ffd6ffe6ff88ff9d000700020000ffe7ffe00000ffdb0004003cffd9ff9d000effe90027002cffee004a0025002affe900130000ffb800890035004c0064ffc4000700000000fff60006ffd8ffea00000000001200270000001400620064001b0000, 1024'h003f003700000000ffb2000000230018ffd0000300470014ffb8fff5fff0ffd6ffe5ff90ff9b0004fff60000ffe8ffde0000ffd9fff5003bffd9ff9b000effea00200026ffea004a001c001fffdf00160000ffb30087003c004e0059ffc7ffff00000000fff60009ffd4ffef000000000012002d0000001d0062005800190000, 1024'h003b003700000000ffb50000001c0017ffcdfff7004c0017ffc5ffecfffbffdaffe3ffa3ffa10000ffee0000ffdfffd20000ffdbffec003bffdaffa8000efffd00220015ffe600520019001fffe1001b0000ffb6007a003f00490046ffce000000000000fff6000cffd1fff200000000001100310000001d005d004800180000, 1024'h003a003700000000ffbc0000001f0010ffd8000000350024ffce000dfffeffe0ffe9ff99ffaf000800000000ffe1ffcd0000ffdb000d003effd4ffae000afff400300026ffe2005700320028ffeb001f0000ffbe006d003a0044004dffca000800000000fff50009ffc9ffde000000000011002c0000000d005c0048001a0000, 1024'h0041003800000000ffb800000027000fffd9001400310020ffc40018ffeeffdcffe9ff85ffa8000d00050000ffeaffda0000ffd90018003dffd1ff9c0008ffdc002c003bffe3004f003a0029ffe6001e0000ffb80079003d00480060ffc2000900000000fff40003ffc9ffdb00000000001200250000000a00630054001b0000, 1024'h0042003900000000ffb0000000290012ffd6000500400018ffb00002fff1ffd5ffe4ff85ff980008ffff0000ffe8ffdf0000ffd90002003cffd7ff97000dffe50027002fffea004c00290029ffe500170000ffb4008d003c004f0066ffc2000600000000fff50004ffd5ffea00000000001200280000001300660064001b0000, 1024'h0041003900000000ffaf000000260014ffd6fffe00430018ffadfffefff5ffd5ffe5ff87ff97000600000000ffe8ffdb0000ffd9fffe003bffd8ff9a000fffeb0029002affe9004f0026002affe600180000ffb6008f003a00500065ffc2000400000000fff50007ffd7ffed000000000012002c0000001500650067001a0000, 1024'h0042003900000000ffb0000000270013ffd6000200420018ffb00000fff3ffd5ffe5ff87ff980007ffff0000ffe7ffdc0000ffd90000003cffd7ff99000effe90028002cffe9004e0027002affe500180000ffb5008d003b004f0064ffc2000500000000fff40006ffd5ffec000000000012002a0000001500650064001b0000, 1024'h0041003900000000ffb0000000280013ffd6000000420019ffb0fffffff4ffd5ffe5ff88ff980007ffff0000ffe7ffdc0000ffd9ffff003dffd8ff9a000effea0029002bffea004e00270029ffe600170000ffb5008d003b004f0064ffc3000500000000fff50006ffd6ffeb000000000012002a0000001500650064001b0000, 1024'h0041003a00000000ffb0000000270013ffd60001003f0019ffb10003fff5ffd6ffe4ff85ff9a000600000000ffe6ffdb0000ffd90003003dffd6ff9a000effea0029002cffea00500027002affe600170000ffb5008c003a00500064ffc2000500000000fff60007ffd3ffe9000000000013002b0000001400660064001a0000, 1024'h0042003b00000000ffaf000000270014ffd400040042001bffb20003fff3ffd5ffe5ff83ff99000800000000ffe7ffda0000ffd70003003fffd5ff98000effe7002a002fffe8005100280029ffe300190000ffb3008d003b00510065ffc0000400000000fff6000affd1ffe8000000000014002d0000001700670063001a0000, 1024'h0042003b00000000ffae000000260011ffd300020047001cffb0fffefff3ffd4ffe3ff87ff96000afffe0000ffe6ffd90000ffd7fffe003dffd7ff98000effe80029002dffe50050002b002bffe4001c0000ffb3008e003d00500065ffc0000700000000fff60008ffd4ffec000000000013002d0000001500660063001a0000, 1024'h0042003a00000000ffaf00000026000fffd500000045001affaefffefff5ffd4ffe1ff88ff960009fffe0000ffe4ffdb0000ffd9fffe003bffd8ff99000effea0027002bffe7004e0029002dffe6001a0000ffb5008e003b004f0065ffc1000900000000fff50006ffd6ffee000000000012002b0000001300650065001b0000, 1024'h0042003900000000ffb0000000270011ffd600010043001affae0000fff5ffd4ffe3ff86ff97000900000000ffe6ffdd0000ffd90000003cffd8ff99000effe80028002dffe9004d0027002bffe500180000ffb6008e0039004f0066ffc1000700000000fff40008ffd6ffec000000000012002b0000001500650066001c0000, 1024'h0042003900000000ffb0000000280012ffd6000100430019ffaffffffff4ffd4ffe4ff87ff970008ffff0000ffe6ffdd0000ffd9ffff003dffd8ff99000effe90028002cffea004d0026002affe500170000ffb5008e003a004f0065ffc2000600000000fff40007ffd6ffec000000000012002a0000001600650065001c0000, 1024'h0040003800000000ffb0000000260012ffd400000047001affaffffafff3ffd5ffe5ff8cff970009fffd0000ffe9ffdd0000ffd9fffa003bffdaff9a000effe90028002affe8004c00280028ffe500190000ffb6008c003c004e0062ffc3000500000000fff50007ffd8ffef000000000012002b0000001500640061001a0000, 1024'h003f003700000000ffb200000024000fffd7fffd00440018ffaffffbfff7ffd6ffe3ff8fff990008fffd0000ffe5ffdd0000ffdbfffb0038ffdaff9e000effee00260026ffe9004b0026002cffe800180000ffb900890039004c005fffc4000800000000fff40005ffd9fff200000000001100290000001200610061001a0000, 1024'h003e003500000000ffb4000000240010ffd6000100450019ffb2fffafff4ffd6ffe5ff91ff9b000afffd0000ffe9ffe00000ffdbfffa0038ffdcff9e000dffe900250029ffe9004700250027ffe500180000ffba00860038004a005effc5000600000000fff40008ffdafff1000000000011002900000015005f005d001a0000, 1024'h003c003400000000ffb600000023000dffd9fffc00420018ffb2fffafff9ffd7ffe3ff95ff9d0009fffd0000ffe5ffe00000ffddfffa0036ffddffa3000dffef00240024ffeb00460023002affe900160000ffbd008300350048005bffc7000900000000fff40006ffdcfff3000000000010002700000012005c005d001a0000, 1024'h003c003300000000ffb800000022000effd90000003e0019ffb6fffffff8ffd8ffe4ff93ffa10008ffff0000ffe7ffe00000ffddffff0036ffdcffa3000dffea00230028ffeb004600220027ffe600160000ffbe007f00330047005bffc7000700000000fff40009ffdaffef000000000010002800000014005b005b001b0000, 1024'h003c003300000000ffb900000021000dffd800000040001affb7fffdfff9ffd8ffe5ff95ffa10009fffe0000ffe7ffe00000ffddfffd0035ffddffa4000effea00230027ffe9004600220027ffe600180000ffbe007e003300450059ffc7000800000000fff4000bffdafff000000000000f002900000014005b0059001c0000, 1024'h003c003200000000ffbb0000001f000cffd8ffff0041001affb9fffbfff9ffd8ffe3ff99ffa20009fffc0000ffe4ffdf0000ffdefffb0035ffdeffa6000effec00200025ffe9004400210027ffe600170000ffc0007b003200440056ffc8000900000000fff20009ffdafff200000000000e00290000001500590056001e0000, 1024'h003a003100000000ffbd00000020000affd9ffff0041001bffbafffafffaffd9ffe5ff9dffa3000cfffc0000ffe6ffe20000ffdffffa0034ffe0ffa8000effec00220024ffea004200220026ffe800170000ffc10078003200410054ffca000a00000000fff3000bffdcfff200000000000e00280000001300580053001e0000, 1024'h0038002f00000000ffbf0000001f0008ffdbffff0040001cffb9fffafffaffdaffe6ffa0ffa5000dfffd0000ffe7ffe40000ffe0fffa0032ffe2ffab000dffec00220024ffea003e00240027ffea00160000ffc500750030003f0052ffca000b00000000fff20008ffdefff500000000000d00240000001000550051001d0000, 1024'h0036002d00000000ffc10000001e0007ffddffff003f0017ffb9fff8fffaffdaffe3ffa3ffa6000efffc0000ffe7ffe90000ffe2fff8002effe4ffad000cffed001d0022ffed0038001f0026ffea00140000ffc70073002d003d0051ffcc000c00000000fff30008ffe2fff800000000000d00230000001000510051001b0000, 1024'h0034002b00000000ffc30000001e0008ffe0fffd003b0016ffbbfff9fffcffdbffe6ffa6ffa9000cfffe0000ffe8ffe90000ffe3fff9002dffe5ffb1000cffef001e0020ffef0037001b0024ffeb00120000ffc90070002a003b004fffcf000a00000000fff30009ffe4fff700000000000c002100000011004d0051001b0000, 1024'h0033002900000000ffc50000001b000affdfffff00380015ffc0fffbfffcffddffe5ffa7ffae000afffe0000ffeaffe90000ffe4fffb002affe5ffb3000affed001b0021ffed0036001b0021ffe900140000ffcc006b00290039004cffd0000900000000fff30009ffe3fff500000000000b002200000010004b004d00190000, 1024'h0033002900000000ffc70000001c000affe3ffff00320014ffc20001fffdffdeffe7ffa6ffb1000a00010000ffe8ffe80000ffe50001002cffe3ffb5000afff0001d0021fff00037001a0023ffec00110000ffcd006900260039004cffd1000900000000fff20009ffe1fff200000000000c002100000010004a004e001a0000, 1024'h0022001b00000000ffc600000016000affc40003007c0019ffc3ffa8ffd9ffdefffdfff0ffa30018ffd40000000bfffa0000ffe3ffa800260002ffb2000affeb00140007ffe70019001d0000ffdd001a0000ffc8005a0048002b0020ffe1fff600000000fff60008ffff002a00000000000f001a00000022003e000d000a0000, 1024'h003c002200000000ffdc0000001b0028ffed0026ffa4000b004d00a8ffd8ffd80023ff7f003a0013003800000024fffd0000ffdd0039fffaffc7ffc8fffdffb9001e0092000c00130011ffccffdb00050000ffbeffdbfffd00370038ffc7ffed0000000000050022ffb3ff5b00000000001000080000005e005b000400000000, 1024'h002c003400000000ffb6000000240014ffee0001fffbffff001600070001ffc30000ffebfff0000100010000000000150000ffdc00030000ffd9ffed000c00000014001400130012ffec0012ffff00000000ff9affd90001004affefffc7001100000000ffef0000fffcffe800000000000f0012000000150070000000020000, 1024'h002d003600000000ffb4000000260012ffee0000fffa00050015000a0004ffc30002ffe9fff0fffe00050000000200110000ffdb00060000ffd9ffec000ffffe001b001700120018fff20014ffff00020000ff99ffd80001004afff0ffc4001200000000fff00003fffdffe500000000000f0010000000140074000100030000, 1024'h002e003800000000ffb30000001d001affdb0005000ffff90023ffef0002ffc1fff3fff6ffedfffcffe90000fff9001a0000ffdaffedffffffd8ffea000f00020004000900120011ffd50006ffec00030000ff8dffd00008004cffd8ffc8000d00000000fff1000cfff4fff2000000000011001d000000230078ffe800030000, 1024'h0023003500000000ffba00000012001cffd5fff200270008003cffd00009ffc600030026fff50002ffdd0000fff400010000ffd9ffce0005ffe10002000f00210013ffee00070019ffddfffcfff2000c0000ff92ffb9000d0042ffb3ffd5000900000000ffef0016fff5fffa00000000001100240000002f006affc200010000, 1024'h0016002f00000000ffc80000000d0004ffdbfff7001600110052ffdb0013ffd3fff70042000a0005ffd60000ffea00040000ffe1ffdffffcffe2001600070024000cffe500040014ffef0006fffe00100000ff9eff9000110030ff9affe0001c00000000fff10003fff4fffc00000000000d00140000000c005dffa2ffff0000, 1024'h001a002e00000000ffd40000000a000cffe7fffcffe80006006a000a001fffd9fff7002a0026fff5ffe50000ffe200000000ffe50007fffbffd30021000700250006ffee000c001dffdb0005fffc000a0000ffa4ff7f0000002cff9bffe2001800000000fff1000affe1ffdd00000000000a0016000000110059ffa700030000, 1024'h0022003300000000ffd4000000180017ffef0018ffd0001d0071003b0009ffd90014000300310005000b0000fffcfff50000ffdb0035000dffca001300040000002700220003002600070000000000100000ffa2ff85fffa0033ffbeffd2001100000000fff10012ffd2ffaf0000000000100019000000140066ffb600060000, 1024'h002b003900000000ffc000000027000bffed0027ffe300150045002cfff3ffce0009fff1000d000f000500000004000e0000ffd7002c0007ffcbfff20004ffe80020002f00050018001a00110002000e0000ff92ffa8000c0041ffdbffc3001c00000000fff0fff7ffe2ffc900000000001200090000ffff0078ffd100040000, 1024'h002e003a00000000ffb0000000280011ffec0007fffbfffe001a0005fffdffc1fffeffeeffee0000fffd0000000000170000ffd90005fffdffd5ffea000ffffd0014001500120014fff50017000100030000ff8dffd10007004dffe9ffc2001700000000fff1fff8fffdffea000000000010000e0000000d007bfff900020000, 1024'h002d003900000000ffaf000000270018ffecfffe0000fffd0014fffdfffeffbf0004ffefffecfffc00000000000400140000ffd9fffd0000ffd9ffec001300030017001000150015ffeb00130001ffff0000ff8fffd800010050ffebffc3000f00000000fff1ffff0002ffed000000000011001400000018007a000000020000, 1024'h002c003900000000ffb0000000270016ffec0000fffffffd0016fffeffffffc00002fff0ffedfffffffe0000000200170000ffd9fffeffffffd8ffed001100030016001000150013ffed00140002ffff0000ff8fffd50002004fffe8ffc3001200000000fff1fffd0000ffed000000000011001200000014007afffc00010000, 1024'h002d003900000000ffb0000000270017ffee0000fffcfffd001800040000ffc00001ffeeffef000000010000000200160000ffd90002ffffffd7ffef000f00030017001300140012ffeb0015000100010000ff90ffd30001004fffeaffc3001200000000fff1fffdffffffea0000000000110012000000140078fffe00000000, 1024'h002e003900000000ffaf000000280016ffec0001fffcffff001a00040001ffc00000ffeeffef000000000000000200170000ffd90000fffdffd7ffec000effff0017001600150012ffed0011fffe00010000ff8effd10002004fffe9ffc3001300000000fff20000ffffffe7000000000011001100000016007afffb00010000, 1024'h002d003900000000ffaf000000260017ffec0000fffffffe0019fffd0003ffc00002fff2ffedfffdffff0000000100150000ffd9fffffffcffd7ffed001100020016001000140016ffec0013ffff00010000ff8dffd20000004fffe5ffc3001300000000fff000010001ffec000000000010001400000015007bfffc00030000, 1024'h002d003900000000ffb0000000260017ffec0002fffffffe0018fffe0000ffc00002fff1ffedfffdffff0000000200150000ffd90002ffffffd7ffed001200010015001000130016ffec0015000000010000ff8effd30001004fffe7ffc3001200000000ffeffffe0000ffed000000000010001500000013007bfffd00040000, 1024'h002e003900000000ffb0000000270017ffec0000fffefffe00170000ffffffc00003ffefffedfffdffff0000000200140000ffd900000000ffd7ffec001200020017001100140016ffee0014000100000000ff8fffd50003004fffe9ffc3001100000000ffeffffdffffffeb000000000010001300000015007bfffd00040000, 1024'h002d003900000000ffb0000000260016ffea00000001ffff0017fffdffffffc00002fff1ffedfffefffd0000000200150000ffd9fffd0000ffd8ffec001200020016001000140015ffed0013000000000000ff8fffd40003004fffe7ffc3001100000000fff0ffffffffffed000000000011001400000016007bfffa00030000, 1024'h002c003800000000ffb1000000240015ffebffff000400000016fff80001ffc10002fff5ffebfffffffd0000000000120000ffd9fffbfffeffd9ffed001200030017000e00120015fff10014000100010000ff91ffd50001004dffe5ffc3001300000000ffee00000001fff00000000000100014000000150078fffa00040000, 1024'h002c003700000000ffb3000000230013ffec00030003fffe0015fffa0001ffc1fffdfff3ffeb0000fffd0000ffff00160000ffdb0000fffeffdaffee001000010012000e00100012ffed0017000000030000ff94ffd60000004bffe8ffc4001500000000ffeeffff0001fff200000000000f0015000000100075fffd00040000, 1024'h002c003500000000ffb4000000230014ffeb0001000700010013fff70000ffc20000fff4ffe90001fffd0000000000130000ffdbfffaffffffdcffeb001000000016001000110012fff10012fffe00010000ff97ffda0001004affe9ffc5001200000000ffec00020001fff100000000000f0013000000160073fffc00060000, 1024'h002a003400000000ffb6000000240010ffeeffff000500000010fff80004ffc3fffdfff5ffe90000fffd0000fffe00160000ffddfffe0000ffddffef001000030014000b00120012ffee0018000100010000ff9affda00010047ffeaffc7001500000000ffedffff0004fff500000000000e00120000000f0070ffff00060000, 1024'h002b003300000000ffb8000000220010ffedffff000200020011fffe0002ffc40000fff1ffecffffffff0000000000130000ffddfffeffffffddffed0012ffff0014001000110013ffef0014ffff00010000ff9cffda00010046ffedffc7001200000000ffee00010001fff000000000000d001200000014006fffff00080000, 1024'h002b003200000000ffba000000200011ffedffff000300000012fffb0003ffc4fffffff3ffecfffffffe0000000000130000ffdefffcfffcffdeffef001300010012000e000f0012ffef0014ffff00030000ff9effda00000044ffebffc7001300000000ffed00020002fff200000000000b001300000013006efffe00090000, 1024'h002a003100000000ffbc0000001e0010ffed00010006ffff0012fff70000ffc4fffffff7ffeb0001fffc0000ffff00150000ffdffffafffdffe0ffef001400010010000c000f000fffed0013ffff00010000ff9fffd9ffff0043ffe9ffc9001200000000ffeb00010002fff500000000000b001300000014006cfffc000c0000, 1024'h0028002f00000000ffbe0000001f0011ffeffffe000500000012fff70004ffc6fffefff9ffec0001fffd0000ffff00140000ffe0fffbfffdffe1fff3001200040014000b0010000efff00013000000010000ffa4ffd9ffff0040ffe8ffca001200000000ffe900010003fff500000000000a0010000000110069fffb000c0000, 1024'h0029002e00000000ffc00000001f0011fff100040002ffff0011fffa0002ffc8fffdfff5ffeb0001ffff0000ffff00140000ffe10001fffeffe0fff00011ffff0013000e000f000efff20013ffff00010000ffa6ffdcfffe003fffecffcb001200000000ffe900020002fff300000000000a00100000000f0066fffe000d0000, 1024'h0028002c00000000ffc00000001d0011ffed0003000b0001000dfff40001ffc9fffcfff6ffe80002fffc0000ffff00140000ffe1fffc0001ffe2ffed0010fffd0011000d000d000efff10012fffb00020000ffa8ffe10000003effedffcc001000000000ffe800030002fff800000000000b0013000000120064fffe000e0000, 1024'h0026002b00000000ffc30000001d000dffeefffd000b0002000cfff30005ffcafffcfff9ffe90002fffa0000fffb00120000ffe3fff80002ffe4fff10010000500110007000e000ffff00014ffff00010000ffacffe30001003bffecffcf001200000000ffea00030002fffa00000000000a0011000000110060fffd000d0000, 1024'h0025002900000000ffc60000001b000effef0000000700020010fff80001ffccfffffff8ffed0002fffc0000fffd00100000ffe3fffb0002ffe4fff1000f00020010000a000c000ffff30011ffff00010000ffafffe100010039ffedffd1001000000000ffea00000000fff5000000000009001000000012005cfffc000c0000, 1024'h0024002900000000ffc70000001c000cfff3fffefffe0001000f00040003ffcefffdfff3fff2000200010000fffe00110000ffe500040001ffe3fff4000d00030012000d000e000efff40015000300010000ffb3ffdf00000038fff2ffd1001100000000ffecfffdfffffff100000000000a000e0000000c005b000000090000, 1024'h0016001b00000000ffc600000019001cffd5001100580006fffeff7dffe1ffde0013003bffc30003ffd40000001000060000ffe3ffa7fffb0001ffcf000cffed001afff7000afffb0022ffe1fff2fff70000ffad00000010002bffc6ffe0ffff00000000ffe10011001d002900000000000f000500000024004fffce00080000, 1024'h003c002200000000ffdc0000001b0028ffed0026ffa4000b004d00a8ffd8ffd80023ff7f003a0013003800000024fffd0000ffdd0039fffaffc7ffc8fffdffb9001e0092000c00130011ffccffdb00050000ffbeffdbfffd00370038ffc7ffed0000000000050022ffb3ff5b00000000001000080000005e005b000400000000, 1024'h002b003300000000ffb6000000230013ffed0000fffe0000001500040000ffc30000ffeefff0000200000000000100150000ffdc00000000ffdaffed000c00000013001300130011ffed0012ffff00000000ff9bffd80001004affeeffc7001100000000ffef0000fffeffeb000000000010001300000016006ffffe00010000, 1024'h002d003500000000ffb5000000260013ffeffffefff700010018000b0008ffc3fffeffeafff2fffe00030000fffe00130000ffdc0006ffffffd7ffef000d00030017001400140016ffeb0015ffff00010000ff99ffd6ffff004affedffc6001400000000fff00003fffcffe500000000000f0010000000140072000000020000, 1024'h0028002d00000000ffb30000000b0022ffc5000a003bfff9002dffbefff3ffc2fff7001fffe80008ffd00000000b001f0000ffd9ffbbfff0ffe6ffea0009fffdfff8fffefffe0000ffd5ffeeffda00160000ff90ffc300170044ffbbffd0000300000000ffed0013fffe000d00000000000f00260000002e006dffc2fffa0000, 1024'h000d002200000000ffcb0000fff00004ffceffcc004f00040044ff860030ffd2ffe4007efff70004ffb40000ffd100010000ffecff90ffe6fff8002600080053fff8ffad00050003ffc9fffffff8000c0000ffb0ff9500000028ff6dffee001f00000000ffe2001a000b003600000000000a0023000000240047ff9000000000, 1024'hffff001400000000fff100000004ffecfffafffd0003002a0063ffe50031ffe80000006b00270017ffed0000ffe500070000fff10003fffafff20041fff900230019ffdf0002000100000011000e000f0000ffd2ff67ffea0005ff83fff1002f00000000ffe000140004000200000000000500070000fff1002bff8d000a0000, 1024'h000a001100000000fff50000000cffe9fff9001cffdc000d0060001d000effe2fff6003500360012ffef0000fff8002f0000fff60019ffefffed002afff6fffcfff00005000affe8ffe700080000000a0000ffceff6ffff70006ffacffef002800000000fff2fff9fff9ffed000000000000fff60000fff1002fffa000020000, 1024'h0013001b00000000ffef00000007000ffffbffedffbbfff5007200320028ffdefff9001a0046fff4fff80000ffe100120000fff4000dffeeffdd003000020029fff6fffc0028fffeffb6ffeeffffffec0000ffc3ff78ffdc001effa8fff2001100000000fff60012ffe2ffc000000000000400080000002c003dffb500040000, 1024'h001b002a00000000ffe2000000150027fff80022ffb2001b008d0053000dffe3001f0002004cfffe001900000006fff60000ffde004c000bffc70020fffefff6002a002e000d0021fff8ffe7fff600070000ffacff6bffe8002cffb4ffdc000100000000fff20024ffcbff940000000000100019000000210058ffaa00050000, 1024'h0027003700000000ffc600000024000effed0031ffd8001a005a0038fff5ffd60010fff6001d000a00080000000900080000ffd7003d0008ffc6fffa0001ffe300220031ffff0021001e000dfffe00160000ff93ff94000d003affcfffc7001900000000fff3fffcffdbffbf000000000012000c0000fffa0074ffc100010000, 1024'h002c003a00000000ffb400000026000fffea000cfff800020022000afffaffc60000fff0fff50004fffc0000ffff00140000ffd90009fffeffd3ffea000dfffa00130019000f0014fffe0016000400040000ff8dffca0007004bffe4ffc3001a00000000fff4fff6fff6ffe5000000000012000f0000000a007bffef00000000, 1024'h002c003800000000ffb000000024001affeb00020003fffb0017fffafffeffc10000fff1ffec0001fffd0000000100160000ffd9fffcffffffd8ffed000d00030013001000120010ffea0012ffff00010000ff90ffd700000050ffe7ffc4001100000000fff1ffffffffffef0000000000120016000000160076fffcfffe0000, 1024'h002b003800000000ffb0000000250016ffed0001fffefffe001a00030003ffc1fffdffefffef000300000000ffff00160000ffda0002fffeffd7ffef000a00050016001200120013ffec0014ffff00030000ff92ffd40001004fffe9ffc5001400000000fff20000fffdffe90000000000120013000000120075fffdfffd0000, 1024'h002c003800000000ffae00000024001affe600050003fffe001ffffe0000ffc1fffefff1ffeffffffffa0000000300160000ffd8fffcfffdffd6ffeb000b00000015001300110015ffe9000cfff600050000ff8effd10007004fffe3ffc5000e00000000fff10004fffaffe90000000000120013000000180078fff4fffd0000, 1024'h002a003900000000ffb0000000210019ffe4fffb0008ffff0025fff30006ffc2fffefffffff1fff9fff30000fffc000e0000ffd9fff30000ffd8fff4000f000e001500040011001affe4000dfff900050000ff8effca0008004cffd6ffc9000e00000000fff10005fffbffef00000000001100160000001b0076ffeaffff0000, 1024'h0028003900000000ffb6000000220013ffebfffffffb0008002a00050006ffc60004fffcfffa0000fffe0000fffe000a0000ffd900050002ffd6fff9000f0009001d000d000e001cfff60013000300070000ff93ffc100040048ffdaffc7001400000000fff20002fff8ffe40000000000110015000000110075ffe900010000, 1024'h002c003900000000ffb5000000240011ffeb000bfff800030025000afffdffc40001fff2fff70002fffe0000000000130000ffd9000affffffd4ffef000efffc00150017000f0015fff70014000000050000ff90ffc60004004affe2ffc3001600000000fff1fffdfff7ffe500000000001100110000000f0078ffee00020000, 1024'h002c003800000000ffb2000000250015ffea000200030000001bfffb0000ffc10000fff5ffee0002fffc0000000000150000ffd9fffcffffffd9ffee000f00010015001100120011ffee0012ffff00020000ff90ffd10001004cffe4ffc4001400000000fff00001ffffffed0000000000110014000000160077fff600020000, 1024'h002b003700000000ffb3000000210012ffeb0000000300010019fff90005ffc2fffcfff7ffed0000fffc0000fffc00130000ffdbfffdfffcffdafff0000f00030013000d00100013ffee0014ffff00030000ff94ffd1ffff004bffe3ffc5001600000000ffef00020000fff000000000000f0015000000120074fff800040000, 1024'h002c003500000000ffb5000000200013ffeb0003000400010019fffd0004ffc2fffdfff4ffee0002fffe0000ffff00140000ffdb0001fffdffd9ffef000f000000120010000e0014ffed0016fffc00060000ff97ffd2ffff0049ffe6ffc4001500000000ffec0004fffffff000000000000f0018000000130073fffa00050000, 1024'h002c003400000000ffb600000023000fffec0001000500040014fffa0003ffc2fffefff5ffeb0004fffe0000fffd00140000ffdcfffdffffffdcffec000fffff0015001100110011fff30015000000010000ff99ffd7fffe0048ffe9ffc5001700000000ffeb00030001fff000000000000f0013000000140072fffb00080000, 1024'h002b003300000000ffb700000024000effed0000000500030010fff90005ffc2fffcfff4ffea0000fffd0000fffc00170000ffddffff0002ffddffee001000000012000d00130011ffec0018ffffffff0000ff9bffd9fffe0047ffeaffc6001600000000ffeb00010003fff500000000000e0012000000120070fffe00090000, 1024'h002b003300000000ffb9000000220010ffecffff000400030012fffb0004ffc3fffffff2ffeb0000fffe0000ffff00130000ffddfffcffffffdeffee001300000014000f00100013ffee0013fffe00020000ff9cffdb00000045ffecffc7001300000000ffee00050001fff000000000000c001300000015006ffffe000a0000, 1024'h002b003200000000ffbb0000001e0011ffec0000000500000014fff90001ffc4fffefff5ffecfffefffc0000fffd00110000ffdefffcffffffdeffef001400020010000c000e0013ffee0014fffe00020000ff9effd900000044ffe9ffc8001200000000ffeb00000000fff300000000000b001400000015006dfffc000c0000, 1024'h0029003000000000ffbd000000200011ffeeffff000600010012fff70000ffc60001fff9ffeb0001fffd0000000100110000ffdffffbffffffe0fff0001400020015000c000f0011fff40013000100020000ffa1ffda00020041ffeaffca001100000000ffea00000003fff400000000000b001200000012006bfffb000d0000, 1024'h0029002e00000000ffbf0000001f000ffff000000002fffe000ffff90001ffc7fffffff6ffecfffffffd0000fffe00150000ffe1fffeffffffe0fff0001200020010000a0010000ffff100160003ffff0000ffa5ffdcffff0040ffebffcb001300000000ffe9fffc0003fff600000000000a00100000000f0068fffe000c0000, 1024'h0029002d00000000ffc00000001d0012fff000000001fffe0010fffe0000ffc70000fff2ffee000000000000000000130000ffe10000ffffffe0fff0001100010011000e000f000fffef0013000000000000ffa8ffdefffe0040ffefffcb000f00000000ffe8ffff0000fff200000000000a00120000001300660001000c0000, 1024'h0029002c00000000ffc00000001c000effed000000080003000dfff60001ffc80000fff7ffea0000fffd0000000100110000ffe1fff9fffdffe3ffed0012fffd0013000d000d0010fff50011fffe00020000ffaaffdf0001003dffedffcb001000000000ffe700030003fff60000000000090011000000130065fffd000d0000, 1024'h0027002a00000000ffc40000001e000afff1fffc000a00010009fff10004ffc9fffefffdffe90000fffb0000fffc00140000ffe4fff80001ffe6fff200120004001000050011000cfff000180003fffe0000ffaeffe0fffe0039ffebffce001400000000ffe6ffff0008ffff000000000009000f000000100060fffe000e0000, 1024'h0024002800000000ffc800000020000cfff4ffff0002ffff000cfff70000ffcb0002fff9ffed0003fffe0000fffe00170000ffe5fffb0002ffe7fff2000f00020010000900140008fff200110006fff90000ffb0ffe2fffc0038ffefffd2001200000000ffeafffe0006fff6000000000009000c00000011005cffff000c0000, 1024'h0024002800000000ffc70000001c0010fff5fffffffafffd000e00040003ffcefffefff1fff2fffe00020000ffff00130000ffe500060000ffe2fff4000d0002000f000c0011000dffed00130002fffd0000ffb3ffe0fffd003afff2ffd2000e00000000ffebfffc0000fff1000000000009000e0000000d005a000400080000, 1024'h0016001b00000000ffc5000000180020ffd40011005800050000ff7dffe0ffdf0015003bffc40000ffd50000001400030000ffe3ffa7fffa0001ffcf000cffed001cfff70008fffe0022ffdefff0fffa0000ffad00000012002bffc6ffe1fffb00000000ffe20013001d002700000000000f000700000025004fffce00060000, 1024'h003c002200000000ffdc0000001b0028ffed0026ffa4000b004d00a8ffd8ffd80023ff7f003a0013003800000024fffd0000ffdd0039fffaffc7ffc8fffdffb9001e0092000c00130011ffccffdb00050000ffbeffdbfffd00370038ffc7ffed0000000000050022ffb3ff5b00000000001000080000005e005b000400000000, 1024'h002b003300000000ffb6000000230012ffed000000000001001300010000ffc40001ffefffee000200000000000000140000ffdcffff0000ffdbffeb000cfffe0014001300130011fff000120000ffff0000ff9bffda00000049ffeeffc7001200000000ffee0000ffffffec000000000010001300000016006fffff00020000, 1024'h002c003400000000ffb6000000240011ffeefffdfffaffff001700080006ffc2fffeffedfff3fffe00000000fffe00160000ffdd00030000ffd9fff1000c00050011000f00140014ffe60017000000010000ff9bffd500000049ffecffc7001400000000fff00000fffeffeb00000000000f0013000000140070ffffffff0000, 1024'h0020002100000000ffb5000000100015ffe00009003e00090000ffb1ffe1ffc9001b0027ffd40015fff500000027000c0000ffdaffc1ffe0fff6ffdc000dffe8001c000efff5ffff002efffd000000150000ffa9ffe4000b003affddffc7000d00000000ffdf00000027001900000000000a0013000000130060ffe8fffb0000, 1024'h0009000700000000ffca0000ffeeffe6ffe5ffe2006fffdbffceff490013ffd0ffce007cffb70003ffb50000ffee003d00000000ff88ffbe00180002000b0023ffc8ffa00003ffceffd2002d000a00050000ffd4ffe2fff80019ffa7ffea003100000000ffccffe50059009d00000000fffa000e0000ffdf002dffe500000000, 1024'h0005fff90000000000020000fff1fff40008ffc6000dfff0000effb70057ffe0ffd9004e0002ffedffe40000ffc2002000000010ffd3ffea000e003b0004004affe2ffac0028ffe5ff9000120004ffde0000000affc7ffb9ffffffaa0004001f00000000ffcb00290022003800000000fff2000d000000180002ffe9001d0000, 1024'h0006fffc0000000000150000000d000700060029ffe2002e0056002d000ffff2001600150033002200190000000b00120000fff80036001afffb0026ffeeffe6002100260002fff3fffdffeafff0000500000005ffa3ffdffff3ffd7fff8000600000000ffdd0031ffeaffc500000000ffff000600000013000affbf00170000, 1024'h0007000700000000fffc0000000effe6fffe000dffe30007003e00330001ffe9fff00019002a0024fff20000ffff00340000fffd000dfffafff60020ffec0005fff8000e000affdfffef00090002000a0000ffedff9c00130000ffd9fffa001b00000000fff8ffe6fff3ffea000000000001ffe80000ffef0018ffbcfff90000, 1024'h000f001200000000fff200000005000cfffcffd9ffb2ffef006b0046002dffe5fff9000f004dfff0fff80000ffe600110000fffafffcffe3ffe1002ffffb0033fffbffff002efffdffb1ffe1fff9ffec0000ffd5ff83ffec0015ffb5fffd00050000000000000012ffdfffb6000000000002fff500000036002bffb9fff70000, 1024'h0015002500000000ffeb0000000f002bfffa001bffa30018009d005e0016ffea00240005005ffff2001c00000008fff00000ffe2004d0004ffc9002dfffdfffe0029002a000f0024ffecffdcfff300070000ffb6ff5effe20022ffaaffe4fffa00000000fff9002dffc8ff8900000000000d001600000029004cffa1fffd0000, 1024'h0023003500000000ffd00000001e0014fff2003dffc90019006e0048fff1ffde0014fff7002d000f000f0000000d00040000ffd8004e0005ffc30003fffcffde0023003afffa001d00250006ffff001a0000ff99ff8300070034ffc9ffca001700000000fff5fffeffd2ffb0000000000012000f0000fff6006cffb6fffd0000, 1024'h002b003700000000ffb600000020000fffea0017fff700000029000efff5ffc9fffdfff2fff9000afffc0000000100160000ffda000ffff9ffd1ffe90005fff3000e001e00090010000400140000000a0000ff91ffc300080049ffe2ffc4001b00000000fff2fff5fff3ffe40000000000130011000000050075ffe9fffb0000, 1024'h002b003500000000ffb0000000230013ffeefffb0000fffe001300010008ffc1fffbfff0ffef000300010000fffc00170000ffdb0001fffeffd7ffef000800060012000f00150011ffe7001a000100000000ff97ffd6fffa004fffeaffc4001700000000ffee00010001fff000000000001400170000001400720002fffb0000, 1024'h002c003300000000ffb0000000260011ffe80003000700070017fffb0001ffc00001fff5ffee0006fffe0000000400180000ffd9fff8fffeffdbffe90007fff9001500170012000efff0000ffffa00030000ff95ffd30000004cffe8ffc4001500000000ffef00070003ffee00000000001300120000001a0072fff6fffc0000, 1024'h0025003100000000ffb30000001e000fffdefff6001bfffc001effd50009ffc1fff60016ffebfffcffe20000fff7001d0000ffdeffd7fff9ffe3fff4000c00100002fff500160009ffd4000afff6ffff0000ff91ffc800050046ffc8ffd1001500000000fff100050009000800000000001000130000001e006dffdffffd0000, 1024'h001e003100000000ffc20000001d000bfffaffe9ffec000b002b000b001fffcc000200090007fffe00080000fff200070000ffe1000bfffdffdc0011000d001d001effff00150018ffec001b0011ffff0000ffa6ffb5ffee003effd2ffd0001d00000000fff200040001ffe500000000000d00120000000b0063ffee00020000, 1024'h002d003300000000ffbf000000260013fff20025ffe1000400320028fff4ffca0006ffe300060007000c0000000b001c0000ffdb0028fffcffd0ffeb0006ffe000120032000e000cfffe000cfff900060000ff96ffbbfffc0043ffebffc3001500000000fff10000fff0ffd1000000000010000c0000000b0072ffed00030000, 1024'h002b003500000000ffb2000000250014ffedffff0003fffe0010fff90001ffc00000fff1ffea000100000000000200190000ffdbfffbfffcffdcffeb0010ffff001200110015000fffec00130000fffe0000ff94ffdafffc004dffecffc4001400000000fff000010006fff10000000000100014000000160075000200030000, 1024'h002b003400000000ffb3000000200013ffedfffe0004fffc0010fff80004ffc1fffdfff4ffeafffffffe0000000000170000ffdcfffcfff9ffdbffee00110002000f000c00110011ffe80017ffff00020000ff97ffd8fffd004bffe9ffc5001400000000ffed00000005fff600000000000e0016000000120072000200040000, 1024'h002d003300000000ffb6000000200012ffedfffe0001ffff0014fffd0004ffc1fffffff2ffeefffe00000000fffe00140000ffddfffefffcffdcffee001000010011000f00110012ffeb0015ffff00010000ff9bffd7fffb0048ffeaffc5001400000000ffea00020002fff000000000000d0015000000170071000000070000, 1024'h002d003300000000ffb8000000230011ffed0000000200020014fffb0004ffc2fffffff4ffecfffffffe0000fffd00140000ffddffff0000ffdcffed0011ffff0013000f00140012ffed0014fffffffe0000ff9bffd7fffd0047ffe9ffc6001400000000ffe800030001fff000000000000d0014000000160072fffd000b0000, 1024'h002c003300000000ffb900000024000fffec0000000500050012fff90004ffc30001fff5ffeb0000fffd0000ffff00150000ffddfffd0003ffdeffee0012ffff0015000d00120013ffee0015000000000000ff9cffd800000045ffe9ffc7001400000000ffeb00040002fff200000000000d0014000000140071fffb000a0000, 1024'h002b003200000000ffbb00000020000fffecfffe000500030014fff90004ffc4fffefff7ffec0000fffb0000fffc00120000ffdefffaffffffdefff0001300030012000c00100012ffef0014ffff00010000ff9effd700010044ffe7ffc8001400000000ffeb00010000fff300000000000b001200000014006efff9000c0000, 1024'h0029003100000000ffbd0000001f000fffed0000000500010015fff80002ffc50000fff9ffed0001fffc0000ffff00140000ffdffffbfffeffe0fff1001400020012000b000f0011ffef0013000000020000ff9fffd600000041ffe7ffca001300000000ffec00020002fff300000000000b001300000013006cfff9000c0000, 1024'h0028003000000000ffbf0000001e0010ffef0000000200000014fff90002ffc70000fff8ffeefffffffd0000fffd00120000ffe0fffefffeffe0fff2001300030013000b00100010fff200130002ffff0000ffa3ffd8fffe0040ffe7ffca001200000000ffe9ffff0000fff300000000000a001000000011006afffa000d0000, 1024'h0029002f00000000ffc00000001e0011fff000040002ffff0012fffcffffffc70000fff4ffed0000ffff0000000100130000ffe000020000ffe0fff10012ffff0012000d000e0010fff10014000000020000ffa6ffdb0000003fffedffca001000000000ffe900000001fff300000000000a0013000000100067fffe000b0000, 1024'h002a002e00000000ffc00000001e000ffff000000001ffff0010ffff0000ffc7fffffff2ffed0001ffff0000ffff00120000ffe1ffffffffffe0ffef001100010012000e000f0010fff20014000100010000ffa8ffde0001003ffff0ffcb001100000000ffe9ffff0000fff100000000000a00110000001200660000000b0000, 1024'h002a002c00000000ffc00000001d0012ffee000200060000000ffff60000ffc80001fff6ffe9fffefffd0000000200100000ffe1fffafffcffe2ffed0012fffe0014000d000c0011fff5000ffffd00030000ffa9ffe10003003dffedffcc000e00000000ffe600020002fff4000000000007000f000000120065fffe000e0000, 1024'h0027002b00000000ffc3000000200010fff100000009fffe000afff0ffffffca0001fffbffe7fffcfffb0000000000130000ffe4fffa0003ffe6fff000130004001400050010000ffff200140002fffe0000ffacffe40003003affecffd0000e00000000ffe6fffc0006fffc000000000008000c0000000e0062ffff000f0000, 1024'h0023002900000000ffc6000000220014fff3ffff0004fffb000bfff6fffcffce0003fff7ffeb0001fffc0000000200160000ffe4fffb0006ffe5fff1000e0005001500080015000afff4000f0005fff90000ffafffe60004003affefffd3000b00000000ffeafff90003fff600000000000b000b0000000f005efffe00090000, 1024'h0023002900000000ffc50000001b0011fff4fffefffbfffc000e0005ffffffcf0002fff1fff2fffe00010000000300100000ffe400030000ffe1fff4000d00050012000a000e0011fff10012000300010000ffb2ffe10005003bfff3ffd3000a00000000ffeffffafffffff100000000000a000e0000000c0059000200030000, 1024'h0015001b00000000ffc400000016001fffd3000e005700040001ff7effe1ffe00014003cffc6fffeffd40000001300000000ffe3ffa5fff60000ffcf000cfff0001bfff6000700000024ffdffff1fffb0000ffadffff0013002bffc4ffe1fffc00000000ffe30010001c002700000000000f000500000024004fffcd00030000, 1024'h003c002200000000ffdc0000001a0027ffec0025ffa5000c004d00a7ffd9ffd80022ff80003a0012003700000023fffc0000ffdd0038fffaffc7ffc8fffeffb9001d0091000c00140010ffccffda00050000ffbeffdafffd00370037ffc7ffed0000000000050023ffb3ff5c00000000001000090000005f005b000300010000, 1024'h002b003300000000ffb7000000230012ffed000000000002001400000001ffc40002fff0ffee000100000000000000120000ffdcffff0000ffdbffec000effff0015001200120013fff10012000000000000ff9bffda00000048ffedffc7001200000000ffee0002ffffffec00000000000f001300000016006ffffe00040000, 1024'h002b003300000000ffb700000023000fffedfffeffff0001001400030003ffc3fffefff0fff10000ffff0000fffe00160000ffdd00010002ffdbffef000d00020010000f00130012ffea0018000100000000ff9cffd6ffff0048ffecffc7001500000000ffeffffe0000ffef000000000010001400000014006ffffe00010000, 1024'h002a002e00000000ffb700000019001efff0000d0012ffff0001ffcbfff6ffd00011fffaffcffff100050000fffcffee0000ffdcfff6fff0ffe1ffcd0013ffed0023000f00070024003200030008fff80000ffa10007fff20043ffefffc5001100000000ffd70006000cfff3000000000007001200000014006b001200140000, 1024'h001c001200000000ffbb000000040018ffea0033007bfff2ffa1ff5dffc6ffd5000f0027ff86fffdffee0000003a000d0000ffe7ffdaffed000cffc30017ffcc0009ffe3ffcc000a0040002e0002002c0000ffd0004b001f0027000cffcc000100000000ffbbffe0004e007c00000000fff600250000ffc300430037000d0000, 1024'h0019fff500000000ffde0000ffecffe0ffebffc20077ffc6ff7dff6c000cffd0ffb70034ff98fffeffb40000ffeb004400000015ff7bffdc0028fff1000f003bffbaff980001ffcfffac00440006000300000018004c0020000d0003fff9001700000000ffc5ffcd004c00ac00000000ffea00070000ffe1000a0035000a0000, 1024'h000dffe90000000000130000fff80002000dffa7fffbfffa0002fff8004fffeaffea0015000d0007fffe0000ffca000d00000014ffc3fffd00100025fff70051000bffdc0037ffe5ffaffff00001ffce00000037fff8ffc6fff9ffe4000c000500000000ffc900370003fff500000000fff8fffb0000004fffeeffff001e0000, 1024'h0001fff300000000001500000010fffd000a0034ffe100350046003b000ffffc000a0008002f002e001f0000000b00190000fffa004a0020fff7001affdaffd3002600350002ffee0013fff1ffec000600000015ffb0ffe4ffefffeafff9000a00000000ffd9002dffe8ffc6000000000007fffd00000002fffbffc700100000, 1024'h0007fffe00000000fffb0000000fffd4fffc0004fff20018001d0031000bffe9ffee000d001f0023fff90000000200300000ffff0007fffdfffe0016ffe9fffafff800120003ffe4fff20016fffc00120000ffffffba0012fff9fff3fff7002000000000fffcfff30000fffb000000000001ffe60000fff00008ffd3fff40000, 1024'h000e000a00000000fffb00000004fff8fffcffccffb9fff0005600420034ffe1ffea00090048fff5fff40000ffd8001c00000001ffebffe3ffed002cfffd0035ffe4fffc0033ffeeff9fffe9fffaffe30000ffe2ff96ffe0000effc5000100130000000000080012ffe9ffc300000000fffffff10000003f001cffc9fffb0000, 1024'h0010001e00000000fff6000000040030fffc0010ff9b000e00a60064001cffeb001d0003006bfff4001d0000fffdfff10000ffe700480001ffcc0036fffb0009001900270014001affd4ffd1fff0fffe0000ffc0ff5dffd0001fffaaffedfff700000000fffc0034ffc3ff8000000000000c001e0000003c003dffa500000000, 1024'h0020003000000000ffd7000000160016fff40042ffbf0023007e0059fff2ffe5001cfff8003d0012001a00000010fff70000ffd8005f0006ffc00008fff5ffd7002a0044fff2002300320001fffe00200000ffa4ff760000002effc7ffcc001400000000fff00005ffc9ffa000000000001300150000fff80063ffaffffc0000, 1024'h0030003600000000ffb9000000210003ffe9001dffef0006002c001bfffaffcafff7ffedfffe0006fffa0000fff900170000ffdc001cfffcffcdffe60001ffea00070021000900140004001cfffe000b0000ff95ffbd000a0044ffe3ffc3002300000000ffedfff3ffedffe2000000000011000f0000ffff0075ffe6fffe0000, 1024'h002e003400000000ffb3000000150021ffcafff80029fffa002fffc40007ffc1fff80014ffe9ffefffd10000ffed000b0000ffdaffc50003ffddffe7000f0010fffaffef00150019ffc3fff2ffe2fffc0000ff89ffd00009004bffbbffd4000500000000ffea001cfff4fffe0000000000110029000000410074ffd100040000, 1024'h0012002c00000000ffc60000fffc001effb6ffe700590013005fff840014ffd5ffff0074fffafff6ffa90000ffe6ffef0000ffddff97000dffee0017000c003d0003ffb5fffb0021ffccffe5ffe500140000ff97ff9700200030ff69fff1000100000000ffeb0023fff2001e0000000000100036000000370059ff77fffd0000, 1024'h000a002d00000000ffea0000fff9fff6ffeaffe0ffe400200091000e0046ffedffec00580040fff8ffd60000ffb8ffdc0000ffed000e000bffd10050ffff005b0010ffc3fffd0036ffe70019001200160000ffbbff5400080017ff6cfff8002c00000000fff10003ffcaffdb000000000006001a0000fff60041ff7900050000, 1024'h0022002f00000000ffe7000000140013ffeb0043ffb2003600a40077fff9ffec001ffff600560015001600000008ffe70000ffd900630012ffbc0010fff4ffdb0034004fffee00300037ffeffff300260000ffacff5f000b0021ffbbffd4001000000000fff40017ffabff7c00000000001100120000000a005fff8c00050000, 1024'h002b003800000000ffc3000000220004ffe80029ffea001500480025fff5ffd30001fff8000b0010fffa0000fffa000b0000ffd900270005ffcaffef0001ffe9001900290000001a00210014000100120000ff94ffa70013003bffd3ffc6002300000000ffeefff3ffddffcf00000000001100090000fff90075ffc700050000, 1024'h002c003600000000ffb60000001f000fffe9000400040004001bfffc0000ffc4fffffff7ffeefffffffa0000fffd000d0000ffdb0000ffffffd9ffee001000000012000d000a0019fff60016ffff00080000ff97ffd200070047ffe5ffc6001500000000ffedfffefffcfff000000000000d00160000000f0072fff500060000, 1024'h002d003400000000ffb800000020000fffecfffe000100020015ffff0003ffc30000fff3ffeefffefffe0000fffe000f0000ffddfffffffeffdbffee001300030013000d000e0018fff20018000200040000ff9cffd700020046ffeaffc6001500000000ffebffffffffffef00000000000c0015000000120072fffd00080000, 1024'h002d003300000000ffb9000000230010ffed0001000100020013fffefffeffc20003fff3ffedfffffffe0000000100140000ffddfffe0001ffddffed0014ffff0015001000120012fff100140001ffff0000ff9cffd700020046ffebffc6001100000000ffe9fffe0000fff000000000000c0010000000150072fffb000c0000, 1024'h002b003200000000ffba000000230011ffeefffd000300000011fff80003ffc30000fff6ffebfffffffd0000000000150000ffdefffafffeffdffff0001400030015000c00130010fff000140002ffff0000ff9effd900000044ffe9ffc7001300000000ffea00000004fff300000000000b0010000000130070fffc000b0000, 1024'h002a003100000000ffbc000000200010fff000020003ffff0010fff9ffffffc40001fff6ffeb0001ffff0000000100160000ffdffffefffeffe0fff0001400000013000d0010000efff00015000200000000ffa0ffd9fffe0043ffebffc8001200000000ffeaffff0004fff500000000000b001100000011006cfffe000c0000, 1024'h0029002f00000000ffbd000000200011ffef00000005fffe000ffff70002ffc5fffdfff6ffea0001fffd0000000000170000ffe0fffbfffcffe1fff0001200010012000d0011000cffef0013ffff00000000ffa3ffdcffff0041ffebffc9001200000000ffe900000004fff600000000000a000f00000011006afffe000c0000, 1024'h0029002e00000000ffbf0000001f0011fff100000003fffe000ffffa0003ffc6fffdfff5ffeb0001ffff0000000000160000ffe1fffefffeffe1fff2001200020012000c0010000dffec0014ffff00010000ffa6ffdcfffe0040ffedffcb001100000000ffea00020004fff500000000000a00110000001100660000000c0000, 1024'h0029002d00000000ffc00000001e0011fff000010001ffff0012ffff0002ffc7fffefff2ffee000200000000ffff00150000ffe10000fffeffe0fff00010000000120010000f000efff00012fffe00010000ffa7ffdcfffe003fffeeffcb001100000000ffe900010000fff000000000000a0010000000130066ffff000d0000, 1024'h0029002d00000000ffc00000001e0011fff000010001ffff0011ffff0001ffc7fffffff2ffee000100000000000000140000ffe10001ffffffe0fff0001000000012000f000f000ffff00013ffff00010000ffa8ffddffff003fffefffcb001000000000ffe800000000fff100000000000a00110000001200660000000c0000, 1024'h0029002c00000000ffc00000001e0013ffee00020005fffe0011fff6fffdffc70003fff7ffebfffdfffc0000000300110000ffe1fff9fffeffe2ffee001200010013000b000e0011fff3000efffe00010000ffa8ffe00004003effecffcd000c00000000ffe700000002fff4000000000008000e000000140065fffc000c0000, 1024'h0024002b00000000ffc2000000200012ffeffffe0009fffe000dffefffffffcb0000fffeffeafffdfff90000000200130000ffe3fff70003ffe5fff200120007001500040012000efff100110002fffd0000ffabffe00004003cffe8ffd1000c00000000ffe9fffd0005fffb00000000000b000c0000000f0062fff9000a0000, 1024'h0021002900000000ffc50000001f0011fff2fffe0005fffe000efff6fffeffcf0002fffbffef0002fffc0000000000140000ffe3fffb0006ffe4fff4000c0006001500070013000afff500110005fffb0000ffafffdf0001003affeaffd2000d00000000ffecfffb0003fff800000000000e000c00000010005bfff800050000, 1024'h0022002900000000ffc60000001c000dfff4fffffffbfffe001200040002ffcffffffff4fff4000000000000fffd00100000ffe400040000ffe1fff5000a0004000f000b000f000efff10013000300000000ffb0ffde00000039fff0ffd3001000000000fff0fffcfffffff100000000000b000d0000000d0057ffff00030000, 1024'h0014001b00000000ffc500000016001dffd30010005600070002ff7effe2ffe00013003cffc7fffeffd50000001200000000ffe3ffa8fff80001ffd0000bffed0018fff6000600000022ffdffff1fffb0000ffadfffe0010002bffc5ffe2fffe00000000ffe60012001d002600000000000f000800000023004dffce00020000, 1024'h003b002200000000ffdd000000190026ffec0023ffa6000f004f00a6ffdbffd90024ff84003b0012003700000023fff90000ffdd0037fffaffc8ffcbffffffbb0020008f000a00160012ffccffdb00070000ffbfffd7fffe00350034ffc8ffed0000000000050024ffb3ff5c00000000000f00090000005e005a000000020000, 1024'h002b003300000000ffb9000000230010ffee0002fffd0002001600030001ffc50001fff0fff0000100000000ffff00130000ffdd0002ffffffdbffed000efffe0014001300120012fff30013000100000000ff9cffd700000046ffecffc7001400000000ffee0000fffeffeb00000000000e001100000013006ffffc00050000, 1024'h002b003300000000ffb8000000230010ffee000000000001001200000002ffc40000fff0ffee000000000000ffff00150000ffdd00010001ffdcffed000fffff0012001000130012ffed00160001ffff0000ff9cffd9fffe0047ffedffc7001400000000ffee00000001ffef00000000000f001400000014006f000000040000, 1024'h002d003500000000ffb8000000210017ffef0003fffafffc0015fffa0001ffc50004ffecffe9fff100000000fff900060000ffdd0004fffeffd9ffe7001500010015000c00120020fff6000e0000fffb0000ff99ffe5fffe0048ffedffc8000e00000000ffe90002fffcffe800000000000900110000001700710006000e0000, 1024'h002a002c00000000ffb700000012003cffea002a0028ffeffff7ffa7ffd8ffd4001dfff8ffb7ffde000000000014ffdd0000ffdafffbfff6ffe3ffbf001dffe500260003ffee00390046fffcffff00080000ffa5002e00070042fff8ffc7fff600000000ffc9ffff000d000300000000fffe001d00000005006a002000190000, 1024'h0019000800000000ffbb0000fffb0022ffe8002c009affddff7eff4affa5ffda000d002bff710004ffe10000004d000d0000ffecffc6fffa0014ffbe0015ffdf0009ffcfffbc0005004b003d000b00380000ffea0070004600250022ffd6ffeb00000000ffaeffb60053009f00000000fff700250000ffb00032004500030000, 1024'h001affe900000000ffe30000fff0ffd1fffbff98005cffc2ff66ff90001dffdaffb10021ffa2fffcffbf0000ffd5003c00000020ff7affe00026ffeefffe0052ffc7ff99001affccffba004e001dffea0000003a0060001c0007001b0001001c00000000ffbbffba0048009d00000000ffefffef0000ffe9fff7004a00040000, 1024'h0016ffe20000000000170000fffcfffb000cffb4ffeb0010fffc00140057ffedfff6fff80015fffc00100000ffd0000700000012ffe00007000b0015fff00028000cfff50038fff2ffafffecfff3ffcd000000430001ffbafff3fffb0006000200000000ffc30051fffeffe300000000fff700040000005cffe9000f00210000, 1024'h000dfff500000000001a00000011ffec0001002fffef00480035002d001bfffa0008ffff00200023001a0000fff800080000fffc0040002afffd0009ffe4ffca001d0031fffeffff0014fff9ffeb000300000019ffccffdeffeafff5fff6001800000000ffd7003dffe7ffcb00000000000000080000000dffffffd6001f0000, 1024'h0007fffd00000000000400000010ffcefff90008000b0022000a001e0001ffeafff1000e000d0032fff400000000003200000000fffd000f0009000effeffff4fff6000ffffeffe0fffa001b0001000f00000006ffd10016fff5fffffff9002300000000fffafff100020008000000000000fff10000ffef0006ffdb00000000, 1024'h000900040000000000010000ffffffe90002ffbeffc0ffed004200440033ffe4ffe5000b00420005fff20000ffd4002300000007ffdfffdefff5002efff9003fffdffff60032ffe3ffa7fff50007ffe30000fff3ffa2ffe80007ffd20006001b0000000000090000ffefffd000000000fffdffec00000033000fffd4fff70000, 1024'h0012001800000000fffc0000fffa0031fff90007ff90000000af00670028ffed001200020073ffe400130000fff0fff00000ffee003dfff3ffcb0036fff900110006001e001d001affb7ffc3ffe4fff60000ffc8ff5bffcc001affa2fff7fff200000000fffa003dffbcff7b000000000006001c0000004c0033ffa300000000, 1024'h001d002d00000000ffe10000fff70035ffc1003fffeb001d00c6001afffbffe9001500330050fff2ffd900000003ffe50000ffd7001f000fffc2001bfffbfff300090010ffe80035ffe5ffc7ffc7002c0000ff97ff4700180024ff71ffe9ffee00000000ffee0033ffaaffaa00000000000f003900000032005dff5400000000, 1024'h0008002700000000ffdc0000ffed0006ffaffff90050003100a1ff9c0006ffe9001300a90027000eff9d0000ffeeffda0000ffdeff9b0002ffeb00300004003c0013ffbdffde00240011ffe0fff200340000ffa1ff45003f0011ff35fff9000f00000000ffea0011ffdc000d00000000000d00250000001e0050ff1bfff90000, 1024'hffe3000800000000fffe0000ffe1ffdfffd1ffe5004f001d008eff5f0020ffff000000fc00280012ff8d0000ffd5fff70000fffbff82ffdb000c0057fffb005afff7ff85fff4ffee0016fff1001c00150000ffcdff2c001affe8ff070019003400000000ffe1fff10013004f000000000000fffc0000ffeb0018ff09fff80000, 1024'hffdcfffa0000000000280000ffe5ffd2001effe7ffaf00040099001a00510005ffec009b0079fffcffe40000ffcc001d00000014002dffe2fff6009afff2005effdfffa30011ffe7ffba00250030000200000006ff08ffd4ffd9ff4c0021003900000000fff0ffe60002000c00000000fff3fff40000ffbfffecff63fffa0000, 1024'h000c00080000000000210000000900050027002eff39002000bd00dd001f00010025ffe400a8000a004f0000000500020000fff900a0ffe9ffc60044ffeaffde00200067001c0000000dffe0000cfff70000fff3ff2bffb6fff9ffc5ffed001600000000fff8001effb6ff47000000000001ffec000000110021ffa100060000, 1024'h0028002400000000ffe20000001e0022fff90062ffa7000600790064ffe3ffdb0017ffda00410007001e0000001f00270000ffdf0068fffbffc5fff8fff8ffaf0007005d000dfffdfffbffe5ffe200050000ffa5ff7dffe5002cffd8ffcc000500000000ffed0017ffd1ff9b00000000000d000a00000014005fffbf00080000, 1024'h0025003200000000ffbf0000001a0014ffea000000000007002cfff90009ffc700030005fffbfffefffb0000fffc000c0000ffddffffffffffddfffd0011000700130007000d0016ffe9000bfffd00040000ff9cffc0fffa0041ffd4ffcd001100000000ffed000bfffbffea00000000000c001a00000018006bffe700090000, 1024'h0029003300000000ffc00000001f000efff20008fff300060027000e0003ffc90003fff8fffc000100030000fffe000d0000ffde0012ffffffd8fff9000f000100180012000b0017fffc0018000500070000ffa0ffc30000003fffe1ffc8001700000000ffeafffcfff8ffe500000000000b001000000008006dffef00090000, 1024'h002d003300000000ffbb000000250011ffee000cfffb000200180005fffaffc50002ffefffef000100000000000500160000ffdd0007ffffffdbffea0012fff50016001900110010fff80010fffe00010000ff9bffd400040044ffedffc6001100000000ffebfffffffdffe900000000000c000d000000100072fff8000c0000, 1024'h002b003200000000ffb9000000210013ffeefffd0006fffd000dfff50002ffc30000fff4ffe8fffdfffd0000000000150000ffdefffaffffffdfffef001500040013000900110012ffed0016000100000000ff9effde00000045ffebffc7001100000000ffeaffff0005fff700000000000b001300000013006f0001000b0000, 1024'h002b003100000000ffbc0000001f0013ffef00010003fffe0010fffb0000ffc5fffefff2ffea0001ffff0000ffff00120000ffdffffffffeffdeffee001300010013000f000f0010fff10014000000010000ffa1ffdeffff0044ffeeffc8001100000000ffe900000000fff200000000000b001300000012006c0001000d0000, 1024'h002b002f00000000ffbc000000200012ffed000300080000000efff7ffffffc5fffffff3ffe80001fffd0000000100150000ffdffffc0001ffe0ffec0011fffe0013000e000e0010fff10013fffd00020000ffa3ffe000020042ffeeffc9001000000000ffe800010002fff500000000000b001200000013006affff000c0000, 1024'h0029002e00000000ffbe0000001e000fffeffffc0006ffff000dfff90003ffc6fffdfff5ffea0001fffd0000fffd00130000ffe1fffbffffffe1fff0001100050012000a000f0010fff00016000100010000ffa7ffe000010040ffeeffcb001200000000ffe8fffe0002fff600000000000a00110000001100670001000c0000, 1024'h002a002d00000000ffc00000001f0010fff0000000000000001000000001ffc70000fff1ffee000000000000000000130000ffe100000000ffe0ffef001000000013000f00100010fff10013000000000000ffa9ffde0000003ffff0ffcb001000000000ffe800000000fff000000000000a00100000001300660000000b0000, 1024'h002a002d00000000ffc00000001e0011ffee00000002ffff0012fffd0001ffc7fffffff3ffeefffffffd0000ffff00130000ffe1fffd0000ffe0ffef001000010011000d00100010ffee0011fffe00000000ffa8ffdd0001003fffedffcc000f00000000ffe80001fffffff100000000000a0011000000150066fffd000b0000, 1024'h0027002c00000000ffc10000001e0012ffecffff000900010014fff2ffffffc90003fffdffedfffffff90000000000100000ffe1fff50002ffe3fff0001000040014000800100010fff2000dffffffff0000ffa8ffdc0003003dffe6ffcf000d00000000ffe800020001fff500000000000b0010000000170064fff5000a0000, 1024'h0022002a00000000ffc40000001e000cfff0fffd00090004000ffff10004ffceffff0002ffed0003fffa0000fffe00120000ffe3fff90002ffe5fff5000d0005001500050010000cfff700140005ffff0000ffaeffda00010039ffe5ffd1001300000000ffeafffe0005fffb00000000000c000e0000000b005efff500070000, 1024'h0023002800000000ffc70000001c0007fff4000000020004000bfffc0006ffd0fffcfff8ffef000400000000fffa00130000ffe500020000ffe4fff2000afffe0010000c0010000afff700170004fffe0000ffb3ffdefffa0037ffeeffd0001700000000ffec00000004fff800000000000c000e0000000b0058fffe00070000, 1024'h0024002800000000ffc80000001c0007fff2000200000003000c00030006ffccfffbffeffff1000400010000fffb00170000ffe500040001ffe4fff1000bfffc0009000f0010000bffea0015fffeffff0000ffb2ffe2fff90038fff5ffd0001500000000fff000060001fff400000000000b0012000000110058000400070000, 1024'h0014001b00000000ffc7000000160018ffd4000b005a000afffeff7cffe7ffdd0010003cffc40004ffd50000000b00020000ffe3ffa4fffa0003ffd1000dfff00016fff50009fffd001dffe2fff2fff70000ffae0001000a002bffc7ffe1000300000000ffe50016001e002800000000000f000a00000028004cffd200070000, 1024'h003a002100000000ffde000000180025ffed0021ffa5000b004e00a2ffdeffd90020ff87003a000f003400000020fffb0000ffdf0034fff6ffc9ffcd0000ffbf001c008a000c0014000dffccffdb00050000ffc0ffd7fffd00340031ffcaffee0000000000050023ffb5ff6000000000000d00060000005c0058000000030000, 1024'h002a003200000000ffbb000000210015ffed0003fffd0001001b00030001ffc60002fff1fff3ffff00000000000100120000ffdd00030001ffdbfff0000fffff0014001200110013ffed000ffffd00010000ff9dffd4ffff0045ffe9ffc9000f00000000ffee0004fffcffe900000000000e001400000017006dfff900060000, 1024'h002a003300000000ffba000000220011ffee0001fffe0003001800030002ffc60001fff2fff1000100000000ffff00110000ffdd00030001ffdbfff0000f00010016001100100014fff30014000100020000ff9dffd500010045ffeaffc8001300000000ffee0000fffdffeb00000000000e001200000012006efffa00060000, 1024'h002a003400000000ffb900000027000efff00002fffa00030015000affffffc30003ffeefff2000200020000000400180000ffdd00050002ffdcfff1001100000017001400130011ffef0016000200010000ff9bffd400040046ffefffc7001200000000fff2fffdffffffeb00000000000e000c000000100070fffc00050000, 1024'h0029003300000000ffb70000001e001bffef0003fffdfff50013fff0fff7ffc60008ffefffe9fff300010000fffc00060000ffdcfffcfff9ffdbffe1001400000013000d0015001b000400090006fff40000ff99ffe9fff7004affecffc6000e00000000ffe8fffc0002ffe900000000000d00110000001d0071000600080000, 1024'h0023002600000000ffb50000000a003bfff1002c0035ffe3ffe0ff89ffcdffd800200005ffa9ffdb000100000013ffd80000ffdcfffbfff3ffe7ffb70019ffe2001efff4ffee003500540007000d00000000ffad0042fffb0042fffdffc8fff700000000ffbcfff2001f001f00000000000200250000fffb005e003300130000, 1024'h001e000400000000ffbd0000fffb000dffeb00200091ffe2ff63ff58ffb5ffd800020019ff6ffff0ffe300000041000d0000fff2ffd600060015ffbd0015ffdcfff8ffc2ffc10010002e0055000d00330000fffc0082004300210039ffd8ffef00000000ffabffb4005700ad00000000fff3002b0000ffa90027006300020000, 1024'h0029ffea00000000ffeb0000fff1ffd2fff0ff900052ffd3ff72ffa5001fffd5ffc6000cffabffecffc20000ffd900240000001eff6cffe40028ffe6000d004dffd0ffa60015ffe3ffb800380011ffee0000003f006a0026000000260000000f00000000ffbeffd30037007d00000000ffe2ffee0000000dfffc004700110000, 1024'h0015ffe60000000000200000fffdfffb000dffb7ffed00140005000f004cffedfffc00060015fffe000c0000ffd6000200000013ffdd000b0011001e000200300014fff00033fff4ffbdffecfffcffcf00000042fff5ffc5ffeefff20008000000000000ffc20045fffdffe200000000fff0ffff00000053fff1000000310000, 1024'h0008fff400000000001e00000013fffa00060036fff100330036001c000a0001000a000b0019002600110000fffd00100000fffe00390027fffd0008ffe9ffd00022002b0006fff20022fff0fff2fff900000015ffccffe6ffe8ffeafffb000f00000000ffd1002cffe9ffd2000000000001fffd000000060001ffca00270000, 1024'h0001fff90000000000060000000dffdc0000000a000c001500040012fffcfff1fff5001200080029fff500000002002d000000020006001600080013ffedfffcfff80001fffcffe3fff9001d0005000d0000000cffdd0016fff4ffff0000001700000000fff4ffe800050013000000000000fff40000ffe6fffbffe400000000, 1024'h0004fffb0000000000030000fff7ffe9fff3ffc0ffd8fff0004100340020ffe7ffef001c00420005ffe20000ffea002300000008ffc4ffdeffff002dfff8003cffd9ffee0022ffe2ffa7ffeafffcfff40000fffcffa20006fffeffce0010000a00000000000dfff9fff2ffe200000000fffaffeb000000340003ffc0ffed0000, 1024'hfff1fff800000000000a0000ffdd001cffdeffddffec000000a9ffe70016fff600280089006afff3ffd40000000ffffb0000fffbffa8ffc70002005000000037fff7ffda000fffecffc2ffa3ffeb00040000ffe3ff38fff1fff2ff530019ffea00000000fffb002dfff7ffda00000000fffb000300000054000aff48ffeb0000, 1024'hffd1fff000000000001f0000ffe3fff000130000ffed0014008affae00220016002800d700530002ffe800000002fff80000000affedffc00011006ffffa00310016ffb60000ffdf0035ffee0037000300000000ff23ffd0ffd0ff320019002700000000ffdbfff9002d002000000000fff5ffe50000ffcdfff3ff46fffa0000, 1024'hffd1ffd900000000002b0000fff4ffe10032004afff3fff10019ffa7fff1001b001400930016000bfffe00000020003e0000001a0026ffc500230039fff0ffdbffeeffd60003ffad003c00110033fff200000025ff8fffc7ffc5ff980012002800000000ffcfffd50055005d00000000ffeeffd00000ff8effd3ffb000020000, 1024'hffe6ffd700000000002d0000fff9ffd6004cfff8ffb7ffcdffc900240022ffffffe300090019fff4002400000003005a0000002a0046ffde001d0044fffd000cffc4ffd80027ffb6ffa300400028ffdc00000050ffe7ffb9ffd900180014001700000000ffecffd50046004300000000ffe6ffe00000ffb4ffbc004600020000, 1024'h001efff40000000000220000001400020048ffeeff32ffee001a010b0024ffec000cff5a006afff7007b0000000c00230000000e0094fff3ffe1001bfffeffe500030072003cfff0ffb100000007ffd500000033ffe2ffa900020073ffedfff70000000000060018ffdaff5e00000000fff3ffe900000034fff8006a000d0000, 1024'h0038001600000000ffe4000000220034fff30040ffa7000200440090ffccffd2002dff880036000c003c0000004000210000ffe0003ffffcffd5ffcb0002ff9a00120093001afff7ffefffbcffccfff70000ffc3ffd5ffe900310036ffc9ffdc00000000fffb0032ffceff7000000000000c0009000000640054000600090000, 1024'h0022002b00000000ffc100000017000effecffe2000dfff70013ffdf0013ffc5fff90011ffeefff8ffed0000fff100140000ffe5ffdafff6ffe80000001700200005ffed001b000affd1000e0003fff60000ffa6ffd2fff9003effd3ffd6001200000000ffed0004000c00050000000000080013000000200060fff2000a0000, 1024'h0023002d00000000ffcc0000001a0013fff8ffffffe200040035001a000fffce0005fffa000efffa00090000fff9000a0000ffe3001a0002ffd90009000f000c0015000c00120017ffe700100005ffff0000ffabffb7fff00039ffdaffd2001100000000ffed0007fff4ffd900000000000a0014000000130060ffec000b0000, 1024'h002b003100000000ffc3000000210017ffec001bffee000a0031001bfff5ffcc000affeb0002000600060000000b00100000ffdb00190002ffd5ffee000cffea001b00290009001300030005fff800080000ff9effc20004003fffe7ffc7000c00000000ffec0005ffecffd300000000000d000f00000012006fffe6000b0000, 1024'h002b003300000000ffba0000001f000fffed0002000500000014fff90001ffc5fffdfff7ffeb0000fffb0000fffd00120000ffdefffefffeffddfff0001200030013000b000c0013fff50018000100050000ff9effd700040043ffe7ffc7001500000000ffeafffc0000fff500000000000b00110000000d006efff9000a0000, 1024'h002b003100000000ffbc0000001f0011ffef00010002fffe0012fffe0000ffc4fffefff2ffec0002ffff0000ffff00140000ffdf0000fffeffdeffef001200010012000f000f0010fff00015000000020000ffa1ffdb00000043ffeeffc8001200000000ffe9ffff0000fff100000000000b001300000012006c0000000c0000, 1024'h002b002f00000000ffbc000000210011ffee000000050001000ffff8ffffffc50002fff5ffeafffffffe0000000100120000ffdffffb0000ffe0ffec0012ffff0015000e00110011fff400120000ffff0000ffa3ffde00010042ffedffc9001000000000ffe700000003fff300000000000b001000000015006bfffe000c0000, 1024'h0029002e00000000ffbe00000020000ffff0fffe0004fffe000cfff70002ffc6fffffff6ffeafffefffd0000ffff00150000ffe1fffd0000ffe1fff0001200030011000800110010ffef00170003ffff0000ffa6ffdf00000040ffedffcb001200000000ffe8fffd0005fff800000000000a00110000000f00680001000b0000, 1024'h002a002d00000000ffc00000001e0011fff0ffff0000ffff000fffff0000ffc70001fff1ffeeffff00000000000000120000ffe1ffff0000ffe0ffef001100010012000e00100010fff000130001ffff0000ffa9ffdfffff0040fff0ffcb000f00000000ffe8ffff0000fff100000000000a00110000001400660001000b0000, 1024'h0029002c00000000ffc00000001f000ffff0000000030001000efffdffffffc70002fff4ffed000200000000000300140000ffe1fffdffffffe2ffef0010ffff0014000f000f000efff40013000100010000ffaaffde0001003efff0ffcb001000000000ffe8ffff0003fff300000000000a000f000000120065ffff000a0000, 1024'h0026002a00000000ffc100000020000cfff0fffd000900000009fff00000ffc90000fffdffe90001fffb0000000000160000ffe3fff4fffeffe6ffee001000010012000900140009fff400120003fffb0000ffabffe0ffff003cffebffce001200000000ffe8fffe0009fffc00000000000b000b000000120062fffc000a0000, 1024'h0023002800000000ffc500000018000cffeffffb000afffe000affeb000affccfff8ffffffeafffdfff80000fff900150000ffe5fff6fffcffe6fff400100004000900000011000bffe80013fffffffd0000ffb0ffdffff90039ffe6ffd1001300000000ffe9000500080001000000000009001400000010005bfffd000b0000, 1024'h0026002800000000ffcb0000000f000cffe9ffff000b00050018fff5000dffcefff6fffcfff2fffefff70000fff3000a0000ffe5fffb0000ffe3fff6001000030006000400070013ffe30010fff500060000ffb4ffd9fff90035ffe3ffd2001100000000ffe80011fff9fff8000000000008001e000000190057fff500100000, 1024'h0026002800000000ffd0000000170003ffecffff00080015001e0004000dffcffffbfffcfff8000cfffd0000fff200080000ffe40002000bffe4fff9000c00010013000f00070012fff60014fffc00070000ffb8ffd2fffc0030ffe7ffd1001900000000ffe8000ffff5ffec00000000000a0018000000170057ffed00130000, 1024'h0015001b00000000ffcf0000001a000bffd60013005600140009ff85ffe9ffdf000c0042ffc90010ffd20000000100060000ffe5ffae00010002ffd50009ffed0018fff90008fff9002bffe8fff7fff80000ffb0fff3000d0023ffc1ffe2001000000000ffe100120017002300000000000e00040000001e004cffc200110000, 1024'h0039002000000000ffde000000170024ffed0023ffab000d004a009fffdcffd90020ff8900370012003400000023fffc0000ffdf0034fff8ffcbffceffffffbe001d008900080013000effcfffda00090000ffc3ffd9000000330033ffcaffed0000000000040022ffb7ff6600000000000d0007000000580055000100020000, 1024'h0029003000000000ffbc00000022000fffeffffefffd0001001600040003ffc60000fff2fff2000200000000000000150000ffdffffefffdffdefff0000e0001001400120013000ffff00011000000000000ffa1ffd600000042ffecffca001300000000ffef00010000ffeb00000000000d000e00000015006afffb00050000, 1024'h0029003100000000ffbc000000210012fff00000fffafffe001800030004ffc6fffffff2fff3fffe00000000fffe00150000ffdf0003fffeffdcfff2000f00020011000f00140010ffea00120000fffe0000ff9fffd4fffc0044ffe9ffca001200000000ffee0001ffffffec00000000000d001100000014006bfffc00060000, 1024'h002a003300000000ffbb000000240013ffee0002fffb0005001900070005ffc7ffffffeefff3000000020000ffff00120000ffdd00070004ffdafff0000ffffe0017001500140013ffed0011fffdffff0000ff9dffd4fffd0046ffebffc8001100000000fff00007fffbffe7000000000010001300000016006efffa00070000, 1024'h002b003500000000ffb900000024000affed00000000000a001400060004ffc60001ffedfff0000300020000fff900110000ffdb00060008ffdaffeb0010fffa0015001500130016fff400180001fffe0000ff99ffd6fffc0046ffeeffc5001800000000fff10003fffdffea0000000000120016000000180070fffd00090000, 1024'h002b003500000000ffb90000001b0011ffec00050005fffe000dffe7fffaffc80009ffefffe2ffefffff0000ffeffff90000ffdc00010000ffdbffd90016fff9000d000800100027000c00110009fff40000ff98fff5fff30047fff0ffc5001600000000ffe500000000ffef00000000000c001d0000001c0071000e00100000, 1024'h0028002700000000ffb90000000c002fffef002e0038fff1ffd3ff92ffccffd40026fffbffa3ffdb00030000001cffd60000ffdcfffefff8ffecffb70023ffdb001efff5ffe1003f00540012000e000d0000ffb4004d000a003d000effc6fff800000000ffc0fff1001f002300000000fff800270000ffef005f003e00180000, 1024'h0021000300000000ffc10000fff8000fffe500190096ffd9ff64ff51ffacffd4ffff001dff6cffefffd70000004600100000fff6ffb6fff8001dffbb0022ffe8fff5ffc1ffc20008002c0046000800320000fffe00840051001f0035ffdbffe800000000ffafffb0005600ad00000000ffeb001b0000ffb4002a005700090000, 1024'h001effe900000000fff10000fff9ffe00000ff860049ffc2ff79ff9c001fffd9ffcc001fffadffe6ffc30000ffd9002900000021ff6effea002afff900180066ffdeff950028ffdcffae0034001bffdc0000003b005e0021fffd0016000b000300000000ffbbffc80040008000000000ffe3ffdf0000000dfff80041001e0000, 1024'h000affe30000000000230000000e0008001effc6ffd5000f000600220031fff8001a00000020fffe00210000fff4000600000011fffb001500110021fffe0021002b00000037ffeeffe1ffe80010ffca00000041fff4ffcaffe90000000bfff300000000ffc9002b0006ffd400000000fff4ffee00000040ffee000400290000, 1024'h0005fff300000000001800000013000100070038ffe8001300240013fff30005000d000400140011000600000005001a00000002002f001cfffcfffbffeaffd1000a001f0010ffeb0016ffedfffaffeb0000000effdffff1fff0fff10002000300000000ffdc000cfff0ffe3000000000001fff30000fffe0000ffd800150000, 1024'hfff4fff10000000000030000fffefff4fff3fff80030000cfff8ffd0fff4fffc000b0035fff90011ffe500000015001400000002ffd0000a0017000ffff7000afffdffe1fff8ffedfff9ffff0000000b00000011fff2001dfff2ffe9000efff900000000fff7fff50018002f00000000fffffffd0000fffaffeeffdbfff20000, 1024'hffe1ffe00000000000140000ffedffd8000effcd00160001fff1ffc1000a000d001100620007000affef00000008000100000015ffadffc8002b0020fffd00290003ffd00003ffdb002dfffd002cfffa00000030ffe3ffffffd7ffd2001a001500000000fff8ffe2003b003700000000fff0ffd00000ffeaffd2ffd7ffee0000, 1024'hffe4ffdc00000000002c0000ffedfff2003c0007ffbfffccffecfff400200018ffea001f0011ffda00150000fff0001f000000260034ffcc00130028fffd0009ffd9ffd7001dffd6ffe700140022ffd700000040fff3ffb6ffd7ffef001a001200000000ffe4ffe90030002800000000ffe6ffdc0000ffc2ffc40024000a0000, 1024'hffffffe100000000002400000000002b00300045ffd3fff5ffce0026ffe300190020ffb3fff4ffed005000000032fff70000000c006f00100007ffe6fffdffaf001b0039fff8ffff0025fff5fff7fff3000000460054ffcaffea005bfffdffd500000000ffdb001c000bffe600000000fff400060000ffefffd20065001a0000, 1024'h0018fff300000000000700000009fff8000d00240005ffedff960033ffe1fffbffe1ff8cffc90003001700000010001f0000000b003b00250002ffcdfffeffcdffe90022ffed0001fff0002effea000d0000003200820020fffd0088fff7ffee00000000fff1ffe6fff9001500000000fff400040000ffddffe9007c00140000, 1024'h0034000d00000000fffc0000000dfff9000affb5ffa7fffbffdf00ca0023ffddffe4ff4b001cfffa00340000ffe3fff90000000200300024ffe0fff3000c00230001003d0015002bffa9001dfff0fffc0000001e00470011001c008effedffee0000000000100005ffb8ff9100000000fff80008000000450011007900130000, 1024'h003d002000000000ffdf000000030041ffaa000cfffd001300770044ffd9ffdc001dffbe002b0004ffe50000000fffdd0000ffd8ffc1000dffd4ffc00007ffdc0012005e00020026ffecff88ffa7000c0000ffb1ffd8002f002effeeffe3ffc8000000000000004eff95ff6e00000000000f0022000000ab005bffa7000f0000, 1024'h0007002b00000000ffdd0000ffe6000dffbaffcf004f001c0081ff91002fffe5fff400940013fff3ff9c0000ffc5ffd10000ffe6ff9f0012ffeb00410011006c0005ff91ffeb0036ffd1fff6fff400230000ffacff71002b0019ff460002000b00000000ffea0019ffdc001d0000000000070039000000230044ff53000a0000, 1024'h000a00270000000000010000fff9ffeeffefffffffc6003b00b5004a0031fffa0004004c00640010ffed0000ffccffd10000ffec00370012ffcc0052fff9003a0025fff2ffed0036001d0010001600250000ffccff34000d0003ff75fff5002d00000000fff00004ffb1ffad00000000000600120000fff1003bff5c000b0000, 1024'h0023002a00000000ffec0000001b0002fff8004bffa9002e00910078fff2ffeb0018fff5004d001f001700000005fffb0000ffdf00660006ffc1000afff2ffd1002c0055fff500190048fffb0002001c0000ffb3ff660008001bffc6ffd2002100000000ffee0000ffb8ff8800000000000bfffb0000fff4005bff96000b0000, 1024'h002a003000000000ffc400000021000cfff00026ffeb000400310019fff4ffcefffefff200000007000000000004001a0000ffdf0022fffcffd4ffee0006ffe7000f00240007000d00080011fffc000a0000ff9effbb0007003bffe2ffc9001900000000ffeafff5fff0ffde00000000000b00070000fffc006cffe300090000, 1024'h002a003000000000ffba000000200017ffeffffd0002fffb0011fffb0001ffc50002fff3ffecfffcffff0000000300130000ffdffffdfffeffdefff0001200050015000b00110013ffec0012ffff00010000ffa1ffdd00020044ffecffca000c00000000ffe9ffff0002fff200000000000b001200000014006c000100090000, 1024'h002a003000000000ffbc000000200013ffed0001000300000012fff9ffffffc70003fff5ffecfffdfffd0000000200110000ffdffffcffffffdfffed001200000016000d00100013fff40010000000000000ffa2ffdc00030042ffeaffca000e00000000ffe900000000fff100000000000b001000000013006cfffb000a0000, 1024'h0029002f00000000ffbe0000001f0010fff0ffff00040000000efff90001ffc70001fff6ffebfffdfffe0000000000110000ffe0ffff0001ffe0fff10013000300140009000f0013fff20017000200010000ffa6ffdd00020040ffecffca001000000000ffe8fffd0003fff700000000000a00110000000f0068ffff000b0000, 1024'h002a002e00000000ffc00000001f000ffff000000000fffe000fffffffffffc70000fff1ffed0000ffff0000000000130000ffe1ffffffffffe0ffee001200000011000e00100010fff20014000200000000ffa7ffdf0001003ffff1ffcb001100000000ffeafffe0001fff100000000000a00110000001200670001000b0000, 1024'h002a002d00000000ffc0000000180016ffe5ffff000cfffb0018ffec0001ffc8fffbfffcffecfff8fff00000fff9000f0000ffe1ffef0000ffe0ffed001200050008000300100012ffe30008fff6fffe0000ffa4ffdc00030040ffe0ffd0000a00000000ffe70006fffbfff700000000000a00170000001f0066fff2000d0000, 1024'h0023002c00000000ffc600000009001dffcdfff8002d00000037ffc1000bffcffff50026fff0fff1ffcd0000ffeb00010000ffe1ffcb0008ffe4fffa0012001affffffe20008001bffcdfff4ffe400060000ffa0ffc600100037ffb0ffe0000100000000ffe7001affef000500000000000b002800000031005fffc0000e0000, 1024'h0017002800000000ffda0000ffe7001bffb3ffec0044000e0079ffa50021ffdeffeb0065000dffeeffa30000ffcfffe30000ffe4ffac000affe40020000e0040fff0ffb6ffef002cffbdffe2ffd5001e0000ffa8ff8a00220021ff65fff8000000000000ffe6002affd2000a000000000005003e0000003a004bff6d00100000, 1024'h000b002200000000fffa0000ffcc000effa9ffed0039002c00ceffb80036fff4ffec009d0042fff8ff920000ffb9ffbf0000ffeaffb4000bffdf004c0005005afff6ffa7ffd6003dffd1ffd6ffd400380000ffbbff36002b0001ff21000d000a00000000ffe20038ffacffef0000000000000045000000350036ff1300160000, 1024'h000500200000000000160000ffe9ffe6ffe60007ffd9005e00dc003800400007000900780071001dffe40000ffbfffb60000ffee0036001bffd10064fff6003c0037ffeaffd70042003e0007001100360000ffdeff0f000cffebff4bfffd003500000000ffdc001dffa2ffa8000000000001001c0000fff0002fff2600210000, 1024'h000c001500000000000300000016fff1ffe0006a000800450089fff1ffdc0006001a005800240031ffde0000fffefff80000ffe800210011ffe5fff8ffeaffbf002d0030ffeaffff0086ffe3fffd00160000ffc3ff70001bfff4ff89ffeb002a00000000ffd60005ffd0ffd200000000000cffeb0000ffe5003fff4a001d0000, 1024'h0037001f00000000ffdf000000180028ffed0021ffaa000a004e0099ffdcffdc0023ff8f0038000e003100000022fff90000ffe00031fff9ffcbffcffffeffc3001e0083000a0015000fffcbffdd00060000ffc2ffd900010032002dffcfffeb0000000000040020ffb7ff6500000000000d0006000000580054fffd00010000, 1024'h0027002f00000000ffbd000000200016ffee0003fffc0000001a00030000ffcb0003fff3fff4fffeffff0000000300110000ffdf00030000ffdcfff1000b000100160010000f0013fff3000effff00020000ffa3ffd600040042ffe8ffcd000d00000000ffeefffefffbffea00000000000d000f000000100068fff700020000, 1024'h0028003000000000ffbc000000200013fff00002fffcffff001700070000ffc90002fff1fff3000100010000000400130000ffdf0004fffeffdcfff2000c000200160011000e0012fff20013000000050000ffa3ffd600050042ffecffcb000f00000000ffeffffdfffdffec00000000000d000f0000000e0068fffb00010000, 1024'h002a003100000000ffbb000000230011fff00000fff9ffff0017000a0003ffc7ffffffeefff3000200010000000100170000ffdf0002fffcffdcfff0000c0000001500150013000effee0011ffff00010000ffa0ffd500020043ffedffca001200000000fff0fffffffdffe800000000000d000c00000012006bfffc00030000, 1024'h002b003400000000ffba000000250013fff00001fff80002001900070007ffc60001ffeefff1fffc00020000000000140000ffde0004fffdffdcfff10011ffff0019001400140013ffeb000efffc00000000ff9bffd400000044ffeaffc9001000000000fff10006fffdffe600000000000b000c00000014006ffffc00090000, 1024'h002a003700000000ffba000000250013ffed0005ffff0003001900020001ffc60004ffefffeffffe00000000000200150000ffdc00040002ffddffef0015fffc0018001300120015ffee0010fffd00010000ff96ffd400020044ffe9ffc7001000000000fff30004fffdffe900000000000d0012000000140074fffa000a0000, 1024'h002a003700000000ffba000000170024ffee000d0001fff00017ffe4fff5ffca0008ffefffe0ffebfffd0000fff7fff70000ffdc0002fff8ffd8ffdf001a000200130005000b0029000c00060003fffa0000ff97fff4fffc0049ffe9ffc7000900000000ffe40000fffaffea000000000007001a000000160072000900110000, 1024'h0023002400000000ffb6000000080039ffeb0037004ffff0ffd0ff7fffbdffda0028000aff99ffe3ffff0000002cffd40000ffdafff6fff9ffefffb30023ffd6002afff6ffd7003c0065000d000600180000ffb5004d0018003b0009ffc8ffec00000000ffbbffee0024003000000000fffd00270000ffea005b003300180000, 1024'h0017000200000000ffc40000000efffcfff30007008fffd8ff54ff51ffb4ffd700000027ff6bffecffd30000003b001f0000fffdffb500080024ffc70021fffefffeffafffdaffff00270057001d001e0000ffff0087005600170035ffe5fff000000000ffb8ff9c006300bd00000000ffeffffd0000ffa60023005700090000, 1024'h0017ffef00000000fff600000014ffe70019ff88000effc4ff75ffd4001cffe2ffe1ffedffbfffdbffe90000ffdd00240000001effa0fffc0021fff50018005bfff3ffb30043ffe4ffc000300033ffbc000000370071000b0005003b0009000000000000ffd4ffc00039004d00000000ffeaffcd0000000dfffb006500150000, 1024'h0008ffeb00000000000f0000000e00290009fff2ffeffff9fff9000dfff3fffb002bffea000dfffa001800000024000c00000003fff10016000dfffcfffffff7001e00150026ffebffe5ffcefff8ffd9000000220014ffeafffd00160006ffce00000000ffe400220005ffdf000000000001fffd00000045fff7000b00090000, 1024'hfff3fff100000000000900000002fffa00030005001f0009fff2ffbffffd000e000b0032ffec0006fff10000fffffffd00000006ffe300000012fffcfff3ffff0010ffe90004fff2002dfff70010fff200000015000affffffefffe5000c000600000000ffe9fffd0017002100000000ffffffee0000fff0ffedffe7ffff0000, 1024'hffeeffec0000000000110000fff9fff7001800120013fff9ffc7ffc800090019fff2000effd7ffef00050000fff6fff700000011001800000012fff9fff7fff7ffffffe0fff6000200220019000ffff90000002e003efff1ffe80011000f000800000000ffeafff5001f003500000000fff5fff60000ffc5ffd4002e00060000, 1024'h0003ffeb0000000000140000fff10002000700160005ffeeffc70021fff00009ffecffc0ffecfff7000c00000012000b0000000e002900160007fff3fffbffe9ffe30004ffe40007ffde0018ffe6001800000039004d0018ffee0050000bffe400000000fffcfff6fff9001600000000fff300100000ffe7ffd2004a00010000, 1024'h0019fffb0000000000110000fff1000afff9ffd7ffdafffa0001005300130006fff0ffaa000fffef000c0000ffdbffd0000000090001000cfff1ffe7000000180002001b00030027fff2ffeaffedfff800000027003e000afffd003c0009ffeb00000000fffd0015ffc1ffb200000000fff700050000003efff2002d00130000, 1024'h001400030000000000040000fffd001dffeb00220000002100220037ffe40001001dffd3000f000a00110000001effdc0000fff100250029ffeeffeffffcffdf0024002fffdb002a0021ffeaffe0002500000009000700250001001dfff6ffdb00000000fff0001affcbffc5000000000001001c0000001a000bfff3000c0000, 1024'h001e001400000000fff70000fffdffe7ffe3ffe2ffe7ffff003500540012ffe6ffd8ffe700260005ffd90000ffda000c0000fffdfffa0011ffe20015ffff0031ffe2fff7fffc0015ffbe0018fff000190000ffedffc7003c000cfff2fffe000b000000000005ffe5ffc1ffde00000000fffc00030000000e0020ffd300020000, 1024'h0007000300000000fff50000ffe7001cffb6ffda003700290086ffcfffeeffef003a006f003a001bffc70000001fffdb0000ffe8ff68ffe1000800120005001d00230004fff2fffe0017ff91ffdd001c0000ffd7ff7d002bfffeff7e0004ffe100000000fff90036ffe3ffcf0000000000050008000000790027ff45fff70000, 1024'hffd0fff40000000000150000ffd7ffc7ffffffd20028ffff006bff70003d0003ffed010400320008ffa50000ffd2001b00000014ffa3ffbb001e008300000070ffdeff690001ffcdffed00190037000a0000fff9ff24fff3ffd0ff140025004400000000ffdfffd8003d007600000000ffeeffe60000ffb9ffefff38fffb0000, 1024'hffe6ffee00000000003d0000fffaffda0054fffeff4efffd0081008e004b00080002003a00920001003c0000ffe7002c0000001c008dffd7fff0008bfff10028fff9fffa002bffd4ffd40024003fffe500000029ff27ff99ffd4ffa6000f003600000000ffebffee0003ffc000000000ffedffd90000ffc2ffe3ffbb000a0000, 1024'h0021000900000000000f00000021002500270067ff3efff9008800daffe9ffed0025ff9c007c0004005a0000002b00340000fff300b3fff1ffc40008ffedff9a00090093002bffe6fff1ffd0ffebffe50000ffdeff76ffb70012000bffdbfff800000000fff1001cffc2ff4e000000000003ffec000000200035ffe6000e0000, 1024'h0029002700000000ffc9000000230030fff50028ffd7fffc0032002fffe9ffcd001cffd3000ffffa001c00000026001a0000ffdc002d0003ffd6ffeb000affd50018003b0014000cffe9ffeeffebfffd0000ffa7ffcafff10040fffbffcbfff100000000ffee0015fff1ffc000000000000e0015000000280064fffc00040000, 1024'h0028003100000000ffb9000000200014ffeefffb0000fffb0013fffafffeffc80004fff8ffeffff8fffb00000002000e0000ffdffffafffeffddfff10011000a0015000600100016fff30014000500010000ffa0ffda00080044ffe7ffcc000d00000000ffedfff60001fff400000000000c000d0000000f006bfffa00020000, 1024'h0028002f00000000ffbc0000001f0017ffee00010000fffc0015fffafffdffc90004fff7ffeffffbfffd0000000600100000ffdffffcfffcffdefff0001100020015000c000f0012fff3000e000000020000ffa2ffd900050042ffe8ffcc000b00000000ffecfffd0001fff100000000000b000f000000110069fff900050000, 1024'h0028002f00000000ffbe000000190016ffe800000008fff9001affef0002ffc9fffcfffeffeefff7fff20000fffc00110000ffe1fff4fffdffdffff200120008000b0001000e0013ffe4000cfff900020000ffa1ffd600050040ffddffd0000b00000000ffeb0002fffdfff800000000000a0014000000160067fff100090000, 1024'h0025002e00000000ffc4000000090021ffd1fffb001ffff9003cffd40008ffccfff5001afff7fff2ffd40000ffef00060000ffe0ffd60002ffdffffc00110019fffdffeb00080019ffcafff5ffe400080000ff9dffc1000f003bffb6ffdc000000000000ffe90014ffebfffb00000000000a00260000002f0063ffc6000b0000, 1024'h0017002900000000ffd30000ffef0022ffb2ffef00480009007aff9f0011ffd9fff8006b000cfff2ffa30000ffe0ffeb0000ffe1ff9f0007ffe7001b000e003dfff7ffbcfff50023ffc0ffd8ffd6001b0000ff9eff8700280026ff64fff7fff800000000ffe80026ffda000a0000000000090036000000420052ff6700080000, 1024'hfff7001700000000fff40000ffd7000affacffe1005d002600b8ff760021fff5000400d900320001ff820000ffd7ffd50000ffecff7bfffdfffa0053000300640000ff8dffe0001cffe5ffceffe9002f0000ffbaff310038fff9ff080018000700000000ffe5001effdd0021000000000002002800000028002cfefb00010000, 1024'hffd4fff70000000000210000ffb7ffe8ffbeffea004e002300e0ff670028001100040130005d000fff730000ffdaffe600000004ff77ffd100110089fff60070ffe7ff6cffd1fff5fffbffce0000003b0000ffeafedf0030ffc3fec70038001d00000000ffe00004fff3004200000000fff0000c0000fff3fff4feb4fff90000, 1024'hffbbffd40000000000520000ffa9ffcafffcffe6ffff001a00dfffa800400026000a013c00900016ffa80000ffe3fffc00000022ffb9ffa9002200bdffee0071ffe4ff75ffdeffcc0005ffe70029002c00000034feb3fff4ff96fed00047003200000000ffd3fff10011003d00000000ffdeffe70000ffc2ffbafecafffc0000, 1024'hffd8ffd700000000006f0000ffe4ffc0006b0011ff18000800c600b600640025fffc006c00cc0008003e0000ffd300260000003200b9ffbdfff000baffe1002ffffbfff70024ffc6fff80022004fffea0000005bfecfff89ffa1ff6c0025004e00000000ffcfffe7ffefffa800000000ffdaffb90000ff99ffbeff74001c0000, 1024'h000bffe80000000000330000001f0030001e00a1ff77000a00920078ffc9000c003dffea006c0010004100000049003e0000fffe0093fff7ffe8fffcffe1ff67001800910028ffbd0023ff9affd6ffda0000ffffff6fffb3ffe4ffd9fff4ffe500000000ffd1003affdaff76000000000001ffd800000020000fff9e00210000, 1024'h0031001e00000000ffe1000000160025ffed001affac000a004e0092ffdeffde0023ff99003b000c002d00000021fff80000ffe1002bfff9ffceffd6ffffffcb001c0079000d0014000dffccffe200030000ffc5ffd4000100300026ffd2ffeb000000000007001dffbbff6c00000000000e0006000000560050fff7fffc0000, 1024'h0024002d00000000ffc10000001e0015fff10002fff5fffd00210006fffeffce0007fff9fffcfffbffff00000003000d0000ffe00004ffffffdbfff6000b00050013000c00110013fff2000d000300000000ffa5ffce0002003fffe3ffd1000c00000000fff1fffcfffcffe900000000000e000e000000120061fff1fffd0000, 1024'h0025002e00000000ffbf0000001f0017fff00004fff4fffc00210008ffffffcd0003fff4fffbfffb000000000002000f0000ffe00008ffffffdafff4000900030012000f00100013fff1000d000100010000ffa3ffd100010041ffe6ffd0000d00000000fff1fffcfffaffe600000000000e000f000000100064fff5fffe0000, 1024'h0027002f00000000ffbc00000020001affee0005fff8fffe001f0008fffcffcb0006fff2fff8fffb000000000007000e0000ffde00060001ffd9fff2000b000200160011000e0016fff1000cfffd00040000ffa1ffd300070044ffe8ffce000800000000fff0fffdfff9ffe700000000000e000f000000120067fff5ffff0000, 1024'h0027003100000000ffba000000240017ffed0000fff9ffff001e00070000ffc90003fff4fff6fffbfffd0000000700110000ffde0000ffffffdafff4000f00070019000f00100016ffef000dfffd00050000ff9dffd1000c0044ffe6ffce000a00000000fff4fffdfffbffe800000000000d000900000010006bfff200010000, 1024'h0026003200000000ffba00000024001affee0000fff9ffff001f00050000ffca0003fff5fff6fffcffff0000000700110000ffdd0000fffeffdafff500120006001c001200110013fff2000bfffd00030000ff9affce00070045ffe3ffcc000a00000000fff5fffefffcffe700000000000e000800000012006dfff000050000, 1024'h0025003300000000ffba000000210017fff00002fffafff7001f0005fffaffc80004fff5fff80001ffff0000000200190000ffdd00040000ffdafff5000f00050011000f0012000dffed0012000300000000ff96ffcc00000045ffe4ffcb000f00000000fff4fff5fffeffec000000000011001000000013006dfff500030000, 1024'h0026003300000000ffb9000000160026ffee000c0000fff20017ffd8fff5ffd0000ffff8ffe0ffe3fffe0000fff6ffed0000ffddfffefff2ffdaffd90016fffd00180005000d002a001afffc0006fff30000ff98fff8fff50047ffe3ffcb000700000000ffe00001fffdffe9000000000007001300000018006e000700110000, 1024'h001c002500000000ffb9000000180032ffeb003c0057fffcffc1ff75ffc6ffe10021000cff94ffdefffa0000002cffe10000ffddffff0011fff5ffb80020ffd3002effeeffe30037005400170005000f0000ffb80052001800380007ffccffed00000000ffc6fff50029004200000000000500220000ffdc0058002f00110000, 1024'h0017001000000000ffc900000016fff9ffedfffa0076ffddff70ff81ffcfffdaffe70004ff82fff2ffcc0000001400240000fff9ffc200250012ffd2001a0011fff2ffb6fff00004fff40051000f000e0000ffee0079005000220033ffeafff600000000ffdcffb2003b009500000000fffe00070000ffc40024004b00020000, 1024'h000dfffa00000000ffee00000004fffefff0ff9e003affebffb4ffbc0009fff0fff80006ffccfff7ffdd0000ffe8fff300000007ff7f0000001affe6000c0044000affd2001ffff9fff3fff80012ffde000000140058001a000a00170008fff400000000fff1fff20018002600000000fffeffee0000003a0000002100020000, 1024'hfff4fff100000000000c0000ffff0005000dfff8000e0003fff0ffd6000a000d000a001ffff5fffc00020000fffdfff600000008fff90009000e000afff6000c0011ffe60006fffb0011ffff0010fff20000001e0010fff0fff2fff4000dfffd00000000ffeb00060014001700000000fffffffd0000fff7ffe6000100000000, 1024'hfffcfff300000000000f0000fffefff7000c0019fff70000ffec000d0002000efff1ffedfff9fffd00070000fffb00050000000a0029000c0000fffbfff0ffeefff60001fff7000200060011fffd000300000020001b0001fff200190009000300000000fff7fff8fffc000900000000fffbfffc0000ffddffe4001900000000, 1024'h0004fff20000000000070000fff60001fffe000100080006ffe40018fff200040008ffdcfff90006001000000015fff500000003000200030007ffeefffbffef00050015ffea000a0011fffefff4001300000023002e0011fff600320001ffef00000000fffd0003fffbfff800000000fffa000400000006ffea0023fffc0000, 1024'h0005fff40000000000070000fff6ffe90002ffe4fff8fff3fff000250000fff5fff3fff4000d000afffc0000000300160000000bffeefff30008000bfffe0014ffe8fffcffffffefffe00012000300090000001dffff0012fff600180005000200000000ffffffe70002000a00000000fff7fff500000001fff0000dfff80000, 1024'h0007fff700000000000b0000fff1000efff5ffdeffe4ffed003600060015fffaffff00130026ffedffee0000ffeafffa00000007ffd1ffe4ffff000cffff001ffff1fff7001dfff6ffd6ffccfff3ffe500000005ffd7ffecfffbffd3000efff500000000fff3001affeeffd900000000fff8fff700000043ffffffd400060000, 1024'hfff1fff700000000000f0000ffea000efff100060008000e0059fff30002fffb001a0057003a0005ffeb0000001e00090000fffdfff6000400050046fffd0019fffeffdcffeefff9ffd2ffecfff2001f00000003ff860009ffeeffa50010ffea00000000fff20011fffe000a00000000fffd001800000008fff7ff97fff50000, 1024'hffe7ffe90000000000180000fff4ffdb0013fff1fffe00200029ffcc0006001700270079001a001bffff00000004ffe50000000bffcfffc0001b001bfff8000c002ffff6fffcffe3008affed003bfffb0000001effafffeeffd3ffab000a002b00000000ffe0ffec0028000700000000fff2ffc30000ffe0ffedffa200040000, 1024'hffddffd50000000000200000fff5ffe30037003e000affcbffbbff9afff3000dffeb0053ffdcfff2fffd0000001a0055000000240027ffcf002b001dfffdffddffc8ffc30004ffb0fffa00340020ffef00000037fffaffd0ffd1ffe80011001a00000000ffcfffc80068008e00000000ffe4ffdb0000ff83ffc6001c000c0000, 1024'h0006ffe500000000002b00000006fff30053ffd2ff78ffc8ffc3009c0036fff5ffdfff8b0029ffdf004f0000ffed00370000002600760007ffff003200070021ffda00040038ffe8ff7a003d001affce000000580027ffb6fff2006f000bfffa00000000fff6ffec0009ffe100000000ffe8fff10000fff2ffcc009800150000, 1024'h0038000800000000000500000022003300090021ff66000d0042010affd9ffe40036ff380060000f00670000003c00090000ffeb0071001dffceffd8fff9ffaa002800b60020000bffe7ffbbffd2fff10000fffefff4ffed0020007dffd9ffc500000000000b0035ffa1ff2500000000000a00020000007a002d003200080000, 1024'h0030002b00000000ffc8000000200014ffe90002ffde000c00290042fff3ffd00011ffc6000d000a00100000000a00020000ffdd0004fffdffd6ffdc0007ffeb0020004300120015000cfff0fff6ffff0000ffafffde0009003d0009ffca000400000000fffb000dffddffae00000000000f0005000000380064fff600000000, 1024'h0026003100000000ffbc0000001c0010ffec00030005fffe0018fff50002ffc8fffdfffcfff0fffcfff90000fffd00110000ffdffffdfffeffdefff3000f0004000c0006000e0012ffe90014fffe00030000ff9fffd4ffff0042ffe2ffcc001200000000fff000020001fff800000000000e0015000000110066fff600010000, 1024'h0025002f00000000ffbf00000010001dffd50000001bfff60032ffd60002ffc9fff50012fff2fff5ffd90000fff3000e0000ffdfffd8fffeffe0fff4000e0010fffbfff3000c0012ffcffff7ffe800040000ff98ffca000c003fffc2ffd9000500000000ffef000ffff3fffb00000000000c001f0000002b0064ffd200040000, 1024'h0017002a00000000ffcc0000fff30027ffb9ffed00410000006affa40012ffd6fff4005c0006ffeeffad0000ffe5fff10000ffe1ffa70002ffe60018000d003cfff6ffc0fff90020ffb9ffdeffd800180000ff9dff960021002eff74fff3fff700000000ffec0022ffe2000c00000000000a00340000003c0053ff8000010000, 1024'hfffd001a00000000ffeb0000ffdc0012ffb1ffe60052001d00adff8a001affef000500bd002f0001ff900000ffe0ffdc0000ffe9ff89fffcfff400490001005b0001ff9dffe2001cffe0ffd1ffe6002f0000ffb5ff4000350004ff200010000200000000ffe8001cffdd001700000000000500290000002b0032ff15fffb0000, 1024'hffd7fffb0000000000130000ffccffeaffc8ffea004c002800c2ff6d001d000d0010011a004d0015ff880000ffe7ffe70000ffffff7fffd700110074fff40062ffffff83ffddfff30018ffd4000c002f0000ffe3fefe002bffd0fee7002c001e00000000ffe1fffe0000003c00000000fff9ffff0000fff20000fed4fff40000, 1024'hffb6ffd500000000003f0000ffc2ffddfff2fff8002f000200b0ff4b00230029000c014700570002ff8b0000ffe600090000001fff8effb7002d008fffec0062ffdeff60fff6ffc1000bffd40024000a00000019fef8fffdffa4fed2004e002500000000ffd5ffe9002e006b00000000ffe9ffd80000ffc8ffc0fedafff40000, 1024'hff9bffae0000000000690000ffa7fff4000d000b0021ffe80097ff3c001c004700150147005bffebffa200000000000900000035ffacffad0045009effe8004fffccff53ffeeffb0fffcffc0001d00020000005eff1cffddff80fee9006c000200000000ffcafff20045007f00000000ffd8ffdd0000ffb8ff79ff02fff70000, 1024'hffa0ff9c0000000000900000ffb2ffd800690011ff9ffff2004cfff800300060001c00ba0072ffee00220000000afff40000004c0062ffba003700a5ffe20032fff9ff9dffe5ffca003e001400550004000000c0ff68ffb1ff68ff86005e001200000000ffc2ffd1003c003a00000000ffc8ffc40000ff66ff49ffa500060000, 1024'hfffaffba0000000000800000fffdffdf008f0058fed3ffd000240165000d002efff4ff5e009ffff000940000001b004d000000420145fff9ffe40051ffd8ffbdffdb006b001bffcfffd4003d0021ffe8000000b0ffbdffb0ffa80083001efffd00000000ffdfffc0ffceff7c00000000ffd2ffb40000ff8cff8b006800190000, 1024'h0033ffe100000000001b000000270050fffe0046ff90ffff001d00c4ffa5fffc0051ff44003f000a00590000006c00160000fff800370012fff0ff9ffff1ff6e003200d1002dffe10011ff71ffb3ffd6000000260035fff70002008bffeeff9800000000fff10048ffb8ff38000000000005ffdc0000009d000c002700130000, 1024'h002d001c00000000ffe300000018001ffff00016ffb1000a00460088ffe2ffe10021ffa00036000c002a0000001cfffc0000ffe30027fffbffd2ffd8ffffffcd0019007100100010000bffd1ffe6ffff0000ffc6ffd7ffff002c0024ffd6fff000000000000a0019ffc3ff7700000000000e000300000051004afff9fffd0000, 1024'h001f002b00000000ffc60000001c0010fff3fffefff2fffe001e0008ffffffd20009fff90000fff9000100000001000c0000ffe30005ffffffdffff8000c0005000e000a00130012fff0000d0007fffc0000ffa9ffd0fffd003bffe6ffd5000d00000000fff8fffbfffeffea00000000000e000f00000012005bfff5fffc0000, 1024'h0021002c00000000ffc40000001d0012fff10000fff1fffd0020000bfffdffd00009fff60001fff9000000000003000e0000ffe100060000ffdcfff6000c0003000c000c00140013ffed000d0005fffc0000ffa6ffceffff003effe6ffd3000c00000000fff7fffafffcffe800000000000f001100000014005ffff4fffa0000, 1024'h0022002e00000000ffc10000001e0013ffeffffdfff3fffe00220006fffdffcf000bfffa0000fff7fffe00000002000a0000ffe000000000ffdcfff5000d00060010000a00150015ffef000a0006fffb0000ffa2ffcd00000040ffe2ffd3000b00000000fff7fffcfffcffe70000000000100010000000180062fff0fffa0000, 1024'h0021002f00000000ffc0000000210012fff0fffffff4000200210005ffffffcf000bfffcfffffff8ffff00000004000c0000ffdf00040002ffdcfff8000d00050014000a00140015fff2000e0007fffd0000ffa1ffca00010040ffe0ffd1000d00000000fff7fffbfffeffea000000000010000e000000110064ffeefffa0000, 1024'h0023003100000000ffbf000000220010fff20001fff10000001e0009ffffffce0008fff6fffcfff9000100000002000e0000ffdf0007ffffffdbfff5000f00020013000e00140014fff300100007fffd0000ff9effcd00000041ffe5ffcf001000000000fff9fffafffeffe800000000000f000c0000000f0066fff4fffd0000, 1024'h0024003200000000ffbd000000220015fff00003fff5fffd001c0006fffcffcc0007fff2fff9fff900010000000400100000ffde00060000ffdbfff2001000000011001000140013ffef000e0003fffd0000ff9bffd2ffff0044ffe8ffcd000d00000000fff9fffcfffeffe90000000000100010000000130069fff8fffe0000, 1024'h0024003300000000ffbb0000001f0014ffed0000fffcfffd001afffffffcffca0007fff6fff5fffafffd00000004000f0000ffddfffefffeffdcfff2001300030010000b00110015ffed000e000200000000ff99ffd300030045ffe6ffcd000c00000000fff9fffdffffffee00000000000f001300000014006afff7ffff0000, 1024'h0023003100000000ffbc0000001d0021ffee000b000cfffc000dffd2fffaffd7000afffdffdbffedfffd0000fff9fff20000ffdefff9fffaffdfffda0013fffa001f0008000e0021001c00020006fff50000ff9dfffafff60042ffe3ffcd000d00000000ffe800060003fff200000000000d00100000001200680002000b0000, 1024'h0013002000000000ffbe0000001f0018fff2002e00570005ffbdff8effcfffdf00150012ffa20004fffb0000002a00080000ffe1fff60012fffeffcd0011ffd70024fff8ffeb000f003e0024000a00110000ffbc003600160032000affd0000100000000ffdeffec0033004b00000000000d00170000ffd60049002300040000, 1024'h0009000700000000ffce00000012ffebfff4ffe7006effdfff7dff70ffe8ffe2ffe5001fff8d0002ffd00000000000290000ffffff9ffff7001dffd0000c0010ffecffc20005ffe6000600350017fff70000ffea00670025001a0019fff0001400000000ffeaffc6004d0088000000000000fff30000ffd80019003dfffa0000, 1024'hfffcfff500000000fff50000fffc00010006ffbd002affd9ffb0ffae001cfff5ffe6000fffcdffe5ffea0000ffe5000c0000000fffb8fff8001afffd00070037ffe8ffbc0020fff1ffc2000e000dffdb00000016004bffef0008000d000efffc00000000fff3fff9002f004600000000fffb000100000010ffed003efffd0000, 1024'hfffcfff300000000000d0000fffa000c0007fffbfff60005ffff001400070007000dfff3000dfffa00110000000cfff7000000040011000f0003000bfff8000100080000fffe0009ffeefff9fff900020000001f000afff9fff70010000affeb00000000fffb0013fffcfff400000000ffff000d0000000cffe7000ffff90000, 1024'h0006fffa0000000000090000fffefff700090009ffe5000c0000002a0000000a0004ffe30009000300150000fffdffec00000003001efffcfff9fff2fff5ffef000d001cfff6000e002e00030007000500000017000f0000fff7001bfffd000800000000fff8fffcfff0ffdf00000000fffbfff50000fff6fff7001000010000, 1024'h0009fff900000000fffd0000fffe0004fffe001a000efff8ffe1fffdffe8fffcffffffe8ffeb0001000500000015000b00000001000b00010003ffe7fffdffe1fff7000efff2fffd00070007fff4000b0000000d0025000b00000023fff9fff600000000fff1fff90006001000000000fffc00050000fff5fffd001f00010000, 1024'hfffeffef00000000fffe0000fffcffeffffeffde002bfffdffceffdcfff4fff400090017ffe90010fff600000016001200000007ffc1fff5001dffff00030010fffeffecfffdffe8ffff000a000b00050000001d001c0014fff600120004fffc00000000fff5ffed0026003100000000fff9fff400000004ffef000efff80000, 1024'hfff1ffe50000000000110000fff4ffe90010ffd50005ffe7ffe7ffcb00130003fff70038fffcfff9ffef0000fff1001300000017ffc2ffd3001f000fffff0021ffebffd6001cffd6fff8fffa001affdf00000026fffeffe7ffe7ffe50015001000000000ffedffef002e002c00000000fff1ffdc00000000ffdffffb00010000, 1024'hfff4ffea0000000000210000fff70015002f0012ffc9ffe6fff5fffd001d00160000fff80004ffd300260000fff2fff400000015004afff8000300110000fffb0001ffee00120005fff90001000effdd000000310018ffbbffea0006000ffff800000000ffdc00110010fffc00000000ffeefffc0000ffe6ffd90035001a0000, 1024'h000affef000000000010000000050021000e005b0009000bffc40014ffc20012001fffb1ffd7fffd00320000003ffff10000fffe005d002b0002ffcbfffeffa0001e003affd3001800450005ffe9001a0000002f0067000ffff30065fff4ffd300000000ffdf0005fffafffb00000000fff800110000ffdbffea005200160000, 1024'h0022000300000000fffd00000011ffd70014ffd9ffdcffe9ff9900810002ffe8ffcdff74ffe8000700160000ffef00240000000e00310028fff5ffed00050015ffe500120003000bffc60058000a00080000002e00670033000b0094fff40004000000000007ffc0ffe7fffe00000000fff6fff60000ffe2fffb008500070000, 1024'h003b001200000000ffed0000001c0015fffaffcaff9e000f001200cafffeffdb001bff580034001300430000000cffee0000ffed000b0008ffdbffd10004fff2002e008300250016fff5ffd2ffecffed0000fff8001e0002002a0072ffd9ffe40000000000110026ffb4ff50000000000009fff7000000840036003c00050000, 1024'h002e002800000000ffcc000000150019ffe20012ffec000600370029fffaffd00002ffd9000c0005000200000003000c0000ffdf0005fffbffd7ffe40005ffe500090035000c000effecffecffe200050000ffabffcdffff0039fff1ffcf000400000000fff6001cffdfffc100000000000d001500000038005dffe700060000, 1024'h0021002d00000000ffc60000ffff001fffbffff70039fffb0051ffb30012ffcdffe90039fff9fff3ffb90000ffdf00050000ffe1ffb70002ffe30002000c0025ffeaffd600050016ffb0ffe9ffd5000c0000ff95ffb000100037ff94ffe7000400000000ffee0025ffe7000900000000000d00330000003f005dffa500070000, 1024'h0003001f00000000ffdf0000ffdf0021ffa2ffe4006b0017009fff700018ffe4fffe00af001b0000ff860000ffdcffe30000ffe3ff720006fff5003700020057fff5ff9cffe9001affc1ffc4ffd400260000ffa5ff5e00300015ff29000cfff900000000ffeb002fffdc001d00000000000b003c00000048003dff25fffb0000, 1024'hffd8000300000000000b0000ffccffeaffc8ffdb0050003300c2ff75002a000b000e0114004b001aff8e0000ffdcffd60000fffaff84ffe3000b007afff00074000cff7effd60005001bffe1001200370000ffe0ff04002dffd9feec0029002300000000ffe50001fff8003400000000fffe000b0000fff10003fedeffed0000, 1024'hffc1ffde0000000000340000ffdaffc70013000bfffa001d0092ffac001d0026001700ff005c0020ffce0000fffa000900000018ffe2ffb7001d007dffe000380008ffa8ffeeffc90058fffe0042001600000021ff0bfff3ffafff1f002d004000000000ffd9ffd5002c003b00000000ffefffc60000ff9cffd0ff19ffec0000, 1024'hffbeffbf0000000000420000fff0ffd200530032ffd3ffee0009ffbb0001002b001c009e0027000d001900000027003d0000002c002bffaa0035004dffe5ffe9fffcffd6000eff9a00540012004dffe500000059ff92ffb1ffaaffa50023002e00000000ffcbffca006e005900000000ffe4ffab0000ff7cffa7ffc3fff80000, 1024'hffc1ffa600000000003f0000fff3ffee004900340019ffb7ff88ff6fffd70023000c0063ffd5fff3000a00000046006800000039fff1ffbc005a000ffff0ffcaffc9ffc8001fff79000100010022ffc9000000780032ffb8ffaf00050030fff700000000ffcfffd3009a00a700000000ffe2ffb80000ffa4ff820033fff70000, 1024'hffadff8e0000000000530000ffdcffe4005bffd70034ffb9ff37ff59fff600320015005affbaffea001b0000003900390000004affbcffc1007c001dfffe000affdaff990019ff8f0002000f0040ffc2000000c10093ffb5ff9a003e004affe700000000ffd8ffd400b500c100000000ffd5ffbf0000ffb4ff440083fff60000, 1024'hffd2ff9a0000000000740000ffe6ffd300a3ffeaff5affa3ff4300840024003bffe3ff810009ffc6008600000003002a0000005c00b0ffda00340025fff5fffaffc9fff50029ffc7ffdb005a004fffb6000000f100abff89ffa100ce0038fffa00000000ffe2ffb80052002600000000ffc7ffb80000ff88ff3d0115000e0000, 1024'h0034ffcc000000000046000000120033004d003eff12ffbaffb50186ffc3fffe0010fe910056ffd900a80000005a003b0000001f00f60037ffdfffcafff4ff82ffd700c30024fff9ff75fff2ffc0ffe00000008f009cffddfff40142fffdff8b000000000009000cffaaff4000000000ffebfffb00000047ffb4010700090000, 1024'h003cfffb00000000ffee0000001d0045ffceffd8fff5001affee006cffb7ffec0052ff6100060009002a00000047ffc70000ffe6ffa7001efffbff8a0007ffc60050009500190019002fff7affc7ffe70000000c007d003000200088ffe9ff9c0000000000050046ffbaff5a00000000000efff4000000cf0025002b00020000, 1024'h0029001c00000000ffe50000001a001bfff10016ffb6000d003f007fffe3ffe30022ffa40031000900280000001cfffc0000ffe40026ffffffd6ffda0003ffce001a006a00100012000cffd4ffe8fffe0000ffc7ffdc000100290024ffd8fff000000000000e0019ffc8ff8000000000000d00010000004b0047fffaffff0000, 1024'h001c002b00000000ffca0000001c000dfff4fffcfff3ffff00180009ffffffd60007fff6fffefff9000100000000000a0000ffe400050001ffe1fff800110005000d000a00130012fff0000f0008fffb0000ffabffd6fffe0038ffebffd7000d00000000fffffffafffeffec00000000000e000e000000100057fff9fffe0000, 1024'h001e002c00000000ffc80000001d000ffff20000fff3ffff001b000afffaffd4000bfff4fffffffa000100000003000c0000ffe200040002ffe0fff500100000000d000e00130011fff1000b0006fffb0000ffa7ffd4ffff003affebffd5000b00000000fffffffbfffdffe900000000000f000f00000015005afff6fffd0000, 1024'h001d002d00000000ffc60000001d000dfff1fffbfff70000001a0003fffeffd30009fffbfffdfffafffe00000001000b0000ffe2fffeffffffe1fff700110005000d000900140011fff0000d0008fffb0000ffa5ffd2ffff003bffe6ffd5000e00000000fffffffb0000ffee00000000000f000f00000013005cfff4fffc0000, 1024'h001e002e00000000ffc60000001f000ffff3fffefff2fffe001d00050000ffd30008fff9fffefff8ffff0000ffff000d0000ffe200030000ffdffff800100005000d000900160011ffed000d0008fff90000ffa3ffd0fffc003cffe4ffd5000f00000000fffffffcffffffeb00000000000f000e00000012005dfff4fffc0000, 1024'h001f003000000000ffc40000001e0013fff10002fff100000021000bffffffd20007fff4fffffff8000100000002000b0000ffe000090001ffdcfff800110002000f000e00120015ffec000b0002fffe0000ffa0ffceffff003fffe6ffd3000b000000000000fffffffaffe600000000000f0011000000120060fff4fffe0000, 1024'h0021003200000000ffc10000001f0013ffed0001fff7000100220008fffdffd10008fff5fffdfffafffe00000002000a0000ffde00030002ffdbfff4001200020011000f00110017fff0000b000100000000ff9bffce00030040ffe4ffd1000c000000000000fffffff9ffe60000000000110012000000160065fff0fffe0000, 1024'h0020003200000000ffc00000001f0013ffee0000fffb00000020fffffffcffd00009fffcfff9fffcfffc00000002000a0000ffdefffeffffffddfff6001200050012000b000f0014fff5000c000500010000ff9affcf00040040ffe1ffd1000e00000000fffefffbfffdffec00000000000f0010000000110065ffefffff0000, 1024'h0020003100000000ffc00000001d0015ffef0003fffbfffa001dfffafffcffd10004fffbfff6fff9fffb0000ffff000c0000ffe00000fffdffddfff300100005000d000800100013fff3000d0005fffe0000ff9cffd400000041ffe1ffd2000f00000000fffbfff9fffeffef00000000000f00110000000e0064fff4fffe0000, 1024'h001f002f00000000ffbf0000001e0027fff00013000ffffc0008ffcdfff8ffe00009fffaffd5ffecfffe0000fff8ffee0000ffdf00020002ffdeffd5000ffff400220009000e00230021ffff0003fff20000ffa00006fff60041ffe7ffd2000800000000ffe900080000fff300000000001000120000000d00610007000c0000, 1024'h0010001e00000000ffbf0000001b001dffe8003300690007ffb7ff7effceffe80010000fff980000fff100000026ffff0000ffe1fff0001cfffeffc3000cffd40020fff2ffe300190040001fffff00160000ffbf004b00200030000cffd6fffb00000000ffe3fff3002c005200000000001000200000ffd70041002300000000, 1024'h0006000700000000ffd300000009ffe4ffedffdb0074ffe7ff81ff7efff0ffe7ffdd001bff940004ffc90000fff5001d00000000ff9f0005001affd9000a0020ffe5ffb8fffafff4fff7003e001200030000fff2006800330017001cfff8001200000000fff5ffc6003d0088000000000002ffff0000ffd9000d003afff50000, 1024'hfffefff600000000fffb0000fff8fff70001ffb40016ffebffcbffdb0021fff8ffec0004ffe8ffeffff10000ffe4fffd0000000dffbbfff40014000300040039fff1ffd10017fffbffd20006000cffe80000001a0035fff90002000f000e0000000000000000fffe0019002100000000fffafffc0000001bffec002bfff90000, 1024'h0004fffb00000000000e0000fff4000e00070004ffd7ffff001e0032001000050002ffe50020fff100140000fffbfff10000000300290004fff3000dfffa0000fffe000bffff0012ffe8fff6fff4000100000013fff2ffedfffc00050004fff300000000fffa0017ffe6ffd700000000fffc000f00000010fff4000700010000, 1024'h000c00010000000000010000fff80013ffea00200009000e00240007ffeb0003000dfff900080002fffb0000000bffe80000fff70006000afff5ffecfff9ffe5000a0019ffea0014001bffe4ffe600130000fffcfffa0012fffffff9fffcffef00000000fff10014ffe0ffe1000000000001000f000000160009ffe200050000, 1024'hffffffff00000000fffe0000fffbfffbfff90001002a000dffedffc400010009fffd001fffdefffeffef0000fff1ffe300000001ffee00090007fff3fffe00080012ffe5ffef00130035000b000c00060000000b001e000efff9fff30002000900000000ffe6fffa0006001e00000000fffd00020000ffe9fffefffa000b0000, 1024'hfffcfff20000000000070000fffefff300050015002b0005ffc6ffd7ffec0009ffff0005ffd50007fffc0000000d000200000007000400100011ffeffffcffee0004fff1ffe800000026001d0007000e0000002300390017ffef001f0003ffff00000000ffe9ffea0015003600000000fff9fffd0000ffd3ffe8001e00060000, 1024'h0008fff400000000000e0000fff9ffee0004ffdffff4ffe6ffdd0021000ffffbffdcffd9fffcfff3fff30000ffe6001000000012fff8000800050003ffff0020ffdbffea000afffdffc30015fffbfff800000027002b0012fff6002a0010fffc00000000ffffffebfff5000b00000000fff3fff800000003ffe5002b00040000, 1024'h000ffffe00000000000f0000ffff001e000afff1ffc40012001d0055000a000a001effbe0021fff4003100000000ffc50000fffd0026000cffeffff40001fffd003200340004002a0025ffdafffdfff60000001b0017ffee00000029fffdffe500000000fff70027ffd1ff9700000000fffd000300000036ffff001a00100000, 1024'h001b000f00000000fff60000000f00030001003dffdb000900080065ffe0fff3fffcffb1000d000d001b0000001c00140000fff300640025ffdefff2fff9ffcd00030038ffe6001400030025ffee00240000fff6fff9002200100038ffe4fff800000000fff8ffeaffd7ffdc000000000004000f0000ffdd001d001800030000, 1024'h0032001d00000000ffde000000080007ffdaffd5ffe8fffb0023004d000bffd8ffebffba0012ffffffef0000ffe1fffa0000ffefffda0002ffddffe300060017fff7002400120018ffceffecffe2ffff0000ffd2fff9001e002a0012ffe7fffd000000000005000effc3ffb4000000000005000a00000056003ffffa00070000, 1024'h001c002000000000ffdd0000ffed002effb3ffed002e000e0082ffcf000bffdc000a00430021fff4ffbc0000ffefffe20000ffe1ffa60004ffe6000f000b0029fffcffe4fff70024ffbfffbbffc800180000ffacff94001d0023ff84fff8ffe700000000fff2003cffcbffdb0000000000080037000000690048ff7800070000, 1024'hffef000f00000000fff50000ffdaffffffb7ffe40063002b00a2ff740012fff6001200e1002f0016ff910000ffeeffe20000ffeeff7afff300060052fffe00580007ff98ffdb00090004ffdafffc00330000ffc6ff350034fff4ff170014001000000000ffe6000dfff50030000000000004001f000000140025ff06fff50000, 1024'hffc5ffe50000000000200000ffdeffc10007ffe8002d0026006eff7b00190017001d0112003b0033ffc10000fff9000600000010ffa5ffbb00290072ffe9004c0013ff98ffefffc4006400070050001400000014ff25fffdffbfff220023004700000000ffd8ffd00042005b00000000fff6ffcf0000ffadffe0ff20ffea0000, 1024'hffbfffc300000000003c0000fff9ffb80068001fffbaffe5fff6ffcd001a0022000500970026001100220000000b005000000032003dffa000300056ffe0fffbffefffcd0022ff8f004800370067ffd400000057ff8fff9affb2ffae001d005000000000ffcbffb5007c006200000000ffe5ff9f0000ff64ffabffe0fff60000, 1024'hffe4ffbd00000000003200000011fffe00740048ff9affb8ff870014fff600150002ffcdfff1ffe200660000003500610000002f008bffce0025fffbffebffa1ffdf00200038ff9ffff700200026ffb40000006c004cff7cffd600650008000300000000ffceffe5006e003300000000ffe7ffc30000ffa5ffa800a400070000, 1024'h000cffd4000000000013000000120030003c0030ffdeffbaff530009ffe40008fff9ff64ffafffc700500000002700250000001b005a00110015ffaeffffffa5ffe8002b0024ffeaffd20003ffe8ffc10000005700e1ffb9ffff00ba0000ffc600000000ffda00120032001700000000fff0fffd00000000ffc300ec00190000, 1024'h0008ffdb00000000000000000008002bfff70013007c0000ff31ff96ffbd00160019ff9cff6effef001900000038ffda00000006ffd900400030ff820006ffb200210015ffe50018003ffff2ffdffff6000000530125001cfffa00b20004ffb400000000ffe2001b0029004500000000000000190000001affc900b400120000, 1024'hfff5ffd700000000001400000005ffcc002bffda00670004fee2ffa2fff5002cffe4ffa8ff52fff8001b0000ffe7ffcd00000023fff500330039ff9f0004fff50019ffd9ffe20020007f00640037ffef00000088014d001fffdc00cf000f000900000000ffe5ffc40043008100000000ffeeffe90000ffa2ff9f00f0001b0000, 1024'h0024ffe20000000000230000000affdb0036fffaffc3ffd4ff1600bbfff10008ffbefed9ffb6ffe200520000fff1001000000025008f0051fffeffa90004ffcfffc40039fff70028ffbb006ffff4fff7000000870130001cfff601470002ffe100000000000fffcaffe1fffa00000000ffe9000a0000ffd7ffac014500180000, 1024'h004dfffe00000000fffe000000120019ffe1ffbaffc00015ffb00110ffc8ffe00026fed20016000f005300000032ffd20000fff200010048ffeaff93000fffd4001a00aa0001003cffd8ffd3ffc400080000003a00c2004700220116ffe5ffa200000000002f0025ff91ff43000000000006001a000000b8000800afffff0000, 1024'h0026001100000000ffde000000110003ffceffbe0026001bfff6fff6ffe6ffec0022ffe4ffe90010ffe90000fff9ffc90000ffebff79fff9ffffffb2000d000b002e002d00120015004cffc20002ffeb0000ffdf003a002d001e0017ffecfff80000000000050010ffe3ffc100000000000bffeb000000730037ffeb00010000, 1024'h0024001c00000000ffe80000001b001afff00011ffbb001100400075ffe9ffe80021ffae00300006002300000019fff90000ffe500210003ffd9ffe00006ffd4001d006100110014000bffd3ffe9fffd0000ffc7ffd900030025001bffddfff0000000000013001bffcaff8500000000000d0000000000480044fff200010000, 1024'h0018002b00000000ffd000000019000dfff3fffffff3000000200009fffeffdc0008fffb0002fff8fffd0000fffe00060000ffe500060003ffe1fffd00140007000b0007000f0014fff0000c0006fffe0000ffaaffd000020033ffe4ffdc000b000000000006fffafff9ffec00000000000d000e0000000e0052ffef00010000, 1024'h0019002c00000000ffce0000001a000ffff00000fff4000300220009fffcffdb000afff90002fffafffe0000000100050000ffe300030002ffe1fff900140002000e000d000f0014fff500060004fffe0000ffa7ffd000020035ffe5ffda000a000000000007fffefff8ffe600000000000e000f000000130056ffed00010000, 1024'h0019002d00000000ffcc0000001a000ffff10001fff80000001f0002fffcffda0009fffdfffefffafffc0000000000070000ffe300020001ffe1fffa00140005000d0008000e0013fff4000b0006ffff0000ffa5ffd100020036ffe2ffd9000c000000000005fffbfffbffee00000000000e000f0000000e0057ffee00000000, 1024'h0019002d00000000ffcb0000001a000efff10000fff70000001e0006fffdffd80005fffafffffffdfffd00000000000b0000ffe300030001ffe1fffb00120005000b000a000f0010fff0000c0005ffff0000ffa6ffd000010038ffe5ffd8000d000000000006fffbfffbffed00000000000f00100000000e0057fff0fffe0000, 1024'h001b002e00000000ffc90000001c000efff2fffefff300000021000cffffffd60007fff80001fffdffff00000000000b0000ffe20003ffffffdffffb00120006000e000d00110011ffee000b0004ffff0000ffa3ffcd00010039ffe5ffd7000d000000000006fffdfffaffe800000000000f000d000000120059fff0fffe0000, 1024'h001b002f00000000ffc70000001e0010fff00000fff4000100240007fffeffd50008fffb0001fffbfffe00000002000c0000ffe10001fffeffe0fffa00120003000f000e00120010fff000070003fffe0000ff9fffca0000003affe1ffd6000d000000000006fffefffcffe700000000000f000c00000013005dffecfffe0000, 1024'h001a003000000000ffc60000001b0014fff00002fff7fffb0024fffefffdffd50007fffffffefff9fffb00000001000c0000ffe10000fffcffdffffb00130007000c000700110011ffee00080004fffe0000ff9dffcbffff003cffdcffd6000c000000000004fffdfffdffed00000000000f001000000010005effecfffd0000, 1024'h001a002f00000000ffc50000001b0018fff00004fffafff90025fffefff8ffd500090000fffefffcfffb00000004000c0000ffe000010000ffdefffb000f0008000d0007000f0010ffee0009000400000000ff9effcc0002003dffddffd70009000000000001fff9fffcffee000000000011001200000010005cffecfff90000, 1024'h001a002f00000000ffc30000001d0015ffef0000fff8fffc0024fffdfffcffd700070001fffdfff8fff90000000000080000ffe1fffeffffffdefff8000c00090011000600120013fff400060005fffd0000ff9fffce0005003dffdcffd9000a000000000001fff9fffbffeb000000000011000c0000000f005cffeafff80000, 1024'h0017002a00000000ffc3000000190022ffee001200160002000affc4fff7ffe8000f0009ffdaffeffffc0000ffffffeb0000ffe0fff9fffcffe4ffd9000bfff10023000600080020002efffc0006fff80000ffa7fffefff80038ffdeffd6000a00000000ffef00080007fffa0000000000110011000000080057fffa00010000, 1024'h0008001800000000ffc800000014000dffef002c00660002ffb4ff7affd5ffec00090020ff9e0001ffec0000001e00070000ffe9ffeb00110005ffd0000bffdd0010ffe4ffe6000c00340028000700130000ffc9003f001900260003ffde000500000000ffe8ffeb0036006400000000000d001a0000ffcc0031001ffffc0000, 1024'h0003000200000000ffdf00000000ffe3fff0ffd5005effe5ff93ff900002ffeaffd60018ffa8fffcffcd0000ffec001d00000005ffa7fffb0019ffe6000b0023ffd8ffb80000fff3ffdf0034000bfffe0000fffb0056002100100014fffe001300000000fffaffd60037007800000000fffd00030000ffe400030036fff80000, 1024'h0001fff60000000000040000ffedfffcfffdffbb0005ffeffff2fffd0021fff5fff200040007fff1fff50000ffeafffb0000000bffccfff6000c001600070039ffe9ffd9000d0000ffba0000fffffff700000019000cfff8fffe0002000ffff800000000000200090007000c00000000fff8000b00000029ffeb0014fffc0000, 1024'hfffdfff50000000000120000fff6000500000000ffe800120034001800010007001c0016002a0007000c0000000affed000000010000fff50001000ffff9fffd00120012fffe0000001affe00002000100000010ffd0fff2fff0ffe40006fffb00000000fff50014fff3ffd600000000fffdfffc0000001afff8ffd300010000, 1024'hfffbfff900000000000b0000fffffff500120018ffebfffe0009ffff00050007fffb00150008000000060000fffb000b000000070025fff6fffe000cfff7fff5fffdfffb0001fff5001600110011fffb0000000dffe5ffeefff4ffed0000001300000000ffe9fff00009000a00000000fffafff40000ffd7fffafff600060000, 1024'h0006fff8000000000003000000050009000e001cfffcfffdffe1fffcfff600030004ffe7ffebfffb00160000000c000100000003002000030002ffeafffcffdf000a0012fffeffff00190004fffffffa000000130029fff0fffe0021fff8fffb00000000ffe90006000a000300000000fffcfffe0000fff2fffa0028000b0000, 1024'h0003fff400000000fffc0000fffffffafff300060034fff7ffceffdfffe7fff3fff8fffdffdf000cffed00000018002300000003ffe0000e0013fff2fffffff5ffe9fff3fff5ffecffe0000dffee000d000000110029001efffd001e0002fff100000000fff8fff40015003700000000fffe00070000fffdfff30015fffb0000, 1024'h0005fffd00000000000b0000fff1fff2ffffffadffddffeb00180024003afff8ffdcfffd0021ffedffeb0000ffc2fff80000000fffd7fff4fffc002100000052ffe5ffd900210004ffb2fffc0005ffe600000013ffeefff6fffdffed001500090000000000040003ffe7ffe500000000fff7fff90000002efff3fffb00030000, 1024'h000e000900000000000e0000ffe40035ffd6001affd6000f009c003c000a0002001000070058ffeafff00000fffcffd90000fff100170010ffdb001efff80000fffd0014fff30028ffc7ffb1ffc100160000ffe7ff8e00020002ffaf000affd400000000fffb0047ffa8ff9a0000000000030030000000530012ff9000050000, 1024'h000100110000000000040000ffd70009ffb50001002b002f00b5ffe60008fffe000f007f004e000bffad0000fff1ffd20000ffecffc2000dffeb003ffffb00340000ffd1ffcf0029fff1ffd0ffd900410000ffd4ff4a0042fff3ff560011fff600000000fff7001fffb8ffe6000000000003002c0000002b001dff26fffb0000, 1024'hffe0fffb0000000000190000ffdcffd1ffe4ffde001e003b009dffbf0017000d002200d800530029ffbd0000ffefffdb00000000ffa5ffd6000f0061fff8004f001dffbaffe1fff80054ffeb002d00280000fffaff250020ffcfff34001a002f00000000ffebffeffffe000e00000000fff8ffe80000ffec0000ff11fff70000, 1024'hffcbffda00000000002f0000fff6ffc20042001dffd90006002dffc10009001e001a00b1002f001e00090000000a00250000001d0019ffb100230050ffed0004000cffd4000affb0007600210061ffed0000002fff69ffc1ffbdff840012004c00000000ffceffbe0058004400000000ffedffb20000ff83ffd4ff98fffe0000, 1024'hffe3ffcd00000000002a0000000fffef0071004cffacffbeff96ffeafffb0019fff8fffaffe3ffea004f0000001500510000002b0086ffcb001dffffffedffb3ffe60005002fffa8002800370042ffb7000000530034ff82ffd900380002002400000000ffc1ffcd006c004800000000ffe9ffc30000ff81ffbe008100120000, 1024'h0016ffdf00000000000d00000018002d00400046ffd0ffbbff520029ffe60000ffebff47ffb0ffc9005800000020003300000017008d00270005ffb0fffaff99ffde00320020fff2ffbc0021ffe5ffc80000004e00ddffb8000b00cafff4ffcd00000000ffd5000b0023001500000000fff4000f0000ffeaffd100ff001b0000, 1024'h0036ffff00000000ffef000000100034ffe5fffa0021fff8ff800036ffe2fff2fff8ff34ffaeffdb001d00000009ffda0000fff80010005dfff5ff8f0007ffd200050036fffa0047ffcbfff4ffbafff90000002700f3002b002300c6fff4ffae00000000fff7002dffcbffd400000000000300360000005bfffd00b800160000, 1024'h0027001000000000ffe9000000060006ffc6ffc900480030ffc9001cffeafff8000dffa4ffd00003ffee0000fff9ffae0000ffedffc10052fff8ffba000a0013002b0012ffdc005a0021fffcffe400210000000c0088006800150063fffaffd5000000000009000dffbeffd800000000000900250000004a0013002f00050000, 1024'h000d000900000000fff50000000bffe5ffebffe100380034ffc9ffdafff300150012fff7ffc7000cfff40000ffe7ffab0000fff8ffca00180004ffbe0004000300400009ffe90037009a0009002300040000000c00610037fffd0025fff8001300000000fff6ffedffeffff8000000000004ffed0000fffd000e000b000c0000, 1024'h000d000800000000fffe00000012ffec001a00240006fff6ff8ffff6fffe000effdaffb1ffafffdf000e0000ffddfff5000000090054002ffff7ffcd0009ffe0fff6fff3fff70027001d004e0011fff400000014008800070005005efff6001000000000fff0ffda0004003000000000fff900040000ffaffff9007d001f0000, 1024'h002b000f00000000fff4000000140008fff0fffdfffc000cffad007bffdaffe90004ff4fffe2fffa00240000001dfff60000fff300310051ffefffc60019ffdbffff003effea003affcf001effd8001b0000000c00870041001b00acffeaffcc00000000001d0000ffcdffd2000000000001002900000029000f0084000e0000, 1024'h002d001d00000000ffe600000012fff4ffdeffadfff10019fff4005efff2ffe70016ffa10004000b00050000fff1ffca0000ffedffb9000dffeeffc7001e00190021003b000d002f0023ffeb0008fff90000ffe3003800370021004cffe8fff9000000000021fffaffc8ff9e000000000006fff900000065003a001c00090000, 1024'h000a001500000000ffe3000000070013ffe500020029fffd0009ffb5ffe2fff300190027ffe7fffcffe300000009fff30000ffeeffc3fff6fffeffe50014fffd000afff6000400030023ffe80009fff70000ffc7fff9000b001affd6ffeffffe00000000fffbfffd000b00100000000000080009000000190034ffd900030000, 1024'h001d001a00000000ffec0000001b0016fff3000bffc0000f003e0068ffefffeb001effbc002e0006001d00000015fffd0000ffe800180001ffdfffea0007ffdf001c00540013000e0006ffd5ffedfffb0000ffcaffd60003001f0011ffe3fff30000000000170018ffd1ff9100000000000bfff900000041003cffec00000000, 1024'h0010002800000000ffd700000015000dfff50002fff1ffff00260009fffdffe2000700020008fffafffd0000000200080000ffe80006fffeffe6000500140007000a0007000d000dffef0005000400000000ffafffc80001002cffdfffe2000800000000000efffcfffaffec00000000000c000a0000000a0048ffe7ffff0000, 1024'h0012002900000000ffd500000015000efff30001fff2000000270009ffffffe1000800000007fffbfffd0000000200070000ffe60003fffbffe4000200150005000c000a000d000ffff20003000200010000ffacffc80001002dffdeffdf000900000000000d0000fff9ffe900000000000c000b0000000e004cffe600000000, 1024'h0013002a00000000ffd400000016000efff40003fff4ffff00260005fffdffdf000700020005fffbfffd0000000000070000ffe60005fffeffe4000200150006000a0008000d000efff10007000400000000ffaaffc9fffe002fffdeffde000b00000000000bfffefffbffed00000000000d000d0000000d004dffe800010000, 1024'h0014002a00000000ffd200000019000ffff40003fff4fffe00240006fffcffde0007ffff0003fffefffd00000000000b0000ffe500050000ffe3ffff00120004000a000a000f000cfff100070005fffe0000ffa8ffccffff0031ffe1ffde000c00000000000afffbfffbffeb00000000000e000d0000000d004fffeb00000000, 1024'h0015002b00000000ffcf000000190011fff30002fff2fffe00240009fffdffdd0007fffc0004fffcfffe00000002000a0000ffe50005fffeffe2ffff00100006000c000b000e000efff00006000400000000ffa8ffcd00010034ffe2ffdd000a00000000000bfffcfff9ffe900000000000e000c0000000c0051ffecfffc0000, 1024'h0016002c00000000ffcc0000001a0013fff10004fff6ffff00240006fffdffdc0007fffc0001fffdfffd00000004000b0000ffe30002fffdffe1fffc00100004000f000d000e000ffff10004000000010000ffa5ffcd00030036ffe0ffdb000900000000000afffffff9ffe900000000000f000b0000000e0054ffeafffb0000, 1024'h0015002c00000000ffca000000190013fff10002fffbfffc00230000fffdffdb00040001fffffffffffb00000003000d0000ffe3fffffffcffe2fffe000e0007000d0009000d000cfff00007000100030000ffa4ffcc00030036ffdeffdb000b000000000009fffcfffdffef000000000010000d0000000c0053ffeafff90000, 1024'h0014002b00000000ffca0000001a0012fff20000fff9fffa0024fffefffcffdb000600040001fffefffa00000000000d0000ffe4fffdfffdffe2fffd000b000a000b00060012000bfff000060005fffd0000ffa4ffcc00000037ffdcffdd000c000000000008fffafffeffef000000000012000c0000000f0052ffe9fff60000, 1024'h0012002a00000000ffc90000001c0012fff20000fff8fffe0023fffefffeffdc000900060002fffcfffb00000005000d0000ffe3fffffffeffe2ffff000a0008000e00050012000dffef00060005fffe0000ffa5ffca00020037ffdbffde000a000000000009fffb0000fff0000000000012000b0000000b0051ffe8fff20000, 1024'h0015002a00000000ffc9000000150017fff00003fff8fff90024fff40000ffe000060004fffdfff0fff90000fffd00000000ffe4fffefff7ffe0fff7000b0006000b0002000d0016fff800010002fffe0000ffa6ffd4fffe0036ffd8ffde000a000000000004fffefffdffee00000000000e000d0000000d0050ffecfff60000, 1024'h0011002500000000ffcb000000140022fff0001a001f00020002ffbcfff1ffef000f000dffd5ffeefffc00000004ffe80000ffe4ffff0001ffeaffdb000dffed001f0001ffff0020002dffff0003fffe0000ffb10008fffb0030ffe4ffdd000400000000fff10007000a000700000000000f00150000fffe0049000000040000, 1024'h0005001100000000ffd10000000e0005ffef002100650000ffb0ff84ffd6ffef0008001fffa30003ffe800000020000b0000ffeeffe1000d000bffd7000dffe40008ffdfffe10009002d0029000700190000ffd700400025001b0009ffe6000300000000ffeeffe20036006700000000000600150000ffca0024001ffffc0000, 1024'h0000fffc00000000ffeb0000fff9ffddfffdffc80043ffe2ff9affaf0004ffedffe00015ffbdfffeffdd0000fff100190000000cffadffea001dfff3000f002cffdcffc00001ffeeffe700330019fffd0000000c004900180006001a0001001400000000fffcffcf0037006700000000fff6fff80000ffe4fffa003afff90000, 1024'h0000fff100000000000a0000fffdffff001affd4ffe8ffedffd9000a0015fffd0002ffeefffefff400190000fff900000000000efff4ffed000e0004000600170002fffa001bfff3ffee00020014ffe1000000250024ffdbfffb001f0004fffe00000000fff400030017fffe00000000fff7fff300000014ffec003700050000, 1024'h0009fff800000000000800000003000e000f0020ffdffff2fff90026fff6fffc0001ffd50006fff9001a0000001100140000000300330004fffafff8fffbffddfff7001b0005fff8ffecfffefff3fffa00000010000dffed00000023fffafff200000000fff10008fffdffee00000000fffb00050000fffffffa002400070000, 1024'h0012000200000000fffa0000fff50019ffe2fffd0015fff3000fffee0000fff8fff2fff3fff8ffecffe40000fff1fff40000fffdffe1000afff8ffeb00010005ffedfff800010010ffd5ffe2ffdafffe0000fff80013000d000afff80004ffe800000000fff2001affe4fff600000000ffff001700000032000afff7000a0000, 1024'hfff9fffc0000000000030000ffe3001cffc6fff4006200160033ff890000000c000a005efff3fffaffb90000fff3ffcf0000fff9ff9e0017000d0005fffd00230008ffc3ffe3001b0003ffccffdf00160000fffbffee0028fff3ffa4001affe400000000ffeb0029ffec001f00000000000300260000002ffffaff9900040000, 1024'hffe1fff20000000000230000ffd2ffd7ffe2ffdb0031001a0053ffd100260014ffe70088002f000effaf0000ffd5fff10000000fffc9000f000d005bfff0005cffe2ff96ffda0008ffdc00130005002d00000021ff8b0037ffd1ff820031001100000000fffcffebffe9003a00000000fff7000f0000ffddffd1ff70fff30000, 1024'hffe2ffe100000000003b0000ffccffdbffeaffd8ffe2002500a10025001f001c00130083007d001cffd40000fff1ffe500000011ffc0ffd2000c005bffea003dfff9ffe5ffeeffee000cffc60003001e0000002dff420015ffbcff720031000d000000000004000bffd8ffd100000000fff1ffe60000001effcdff3bffef0000, 1024'hffcbffd40000000000440000ffdeffd0002b0004ffc4001c0074ffff001a0024002a00a9006c001b000a0000001000060000001c000affb5001f006dffee0016000fffe4fffcffc6004afff1003c00050000003eff38ffccffaeff720023002c00000000ffe6fff00029000400000000ffeaffc70000ffc5ffc2ff67fff90000, 1024'hffdaffd00000000000400000000affd400740043ff81ffe4ffed002b000a0020000c00230029000600550000001400440000002a0091ffbc00170031ffedffc7fffe00170025ffa8004b00300054ffcc00000052ffc4ff89ffc200010006003b00000000ffd0ffcb0052001400000000ffe5ffad0000ff7cffc1002800120000, 1024'h000effe10000000000170000001f002300560065ff9dffb3ff83003effdf0003fff3ff65ffd2ffd5006400000024004c0000001900ab00000000ffc1fffaff85ffdf004a0030ffd0ffe00017fffbffb90000003a0090ff9a000200a0ffeeffe800000000ffd3fff9002cfffd00000000fff0ffec0000ffd1ffdf00d300230000, 1024'h0032000100000000ffea0000000c004cfff200170012ffd2ff860022ffdeffe9ffefff3dffaeffcb002100000016fffe0000fff9002e004afff1ff9e000dffc6ffea002a00040030ff9cfff6ffb3fff10000001500db000b002d00b3ffeeffa700000000ffed002cffe0ffec000000000000004300000049000600c300190000, 1024'h0031001600000000ffe20000fffc001dffb6ffc3004b0023ffe8001dfff0ffeb0007ffa6ffddfffaffe00000fff6ffb10000ffe8ffb40055ffeeffc5000d0023001c0008ffde005effe7ffecffcb00260000fffc006f00680022004cfffaffc30000000000050022ffadffd000000000000b003e0000006d001f001c00050000, 1024'h0010001300000000fff20000000cffd8ffd8ffbd002100480025001dfffefffa0021001d00120022ffe10000fff0ffc00000ffefffb30023fffaffff00020037003effffffeb003400570004001d001e0000fff4ffe2005a0000ffebfffe000f000000000009ffe8ffd4ffd6000000000008ffef0000001f0021ffadfff90000, 1024'hfffa000800000000fffc00000019ffd30012fff3ffdc0010000f000b00010002000f002c00130009fffe0000fff8000700000001fffdffe8ffff000b0002000a0016ffff0017fff3004a0016003bffec0000ffeeffc50006fffaffdcfffa002e000000000002ffca0014fffc00000000ffffffc70000ffd40019ffd3fffb0000, 1024'h0001000700000000fff80000001400130021001cffcfffd9ffe9fff7fffbfffe0006ffedfff4ffd50018000000070016000000020034fff0fff7fff70011ffe7fff6ffff0023fff7fff200080012ffd70000ffe8000bffd200100007fff5ffff00000000fffafff2001f000900000000fffcfff20000ffe700130030000a0000, 1024'h000f001200000000ffee00000013002300030016fff0ffeeffe6001fffe8ffee000effbffff2ffe2001600000023000e0000fff400300022fff2fff6001cffeafffd000d00030016ffc3000affec00020000ffe200220008001e0033fff1ffd700000000000f0003fffdfffb000000000002001b00000007001c003c00080000, 1024'h0015001d00000000ffe7000000160008ffecffdcfff6000b0006002afff1ffee0017ffd60002fff8ffff00000007ffe90000ffeeffdf000efff2ffec00210011001d0019000b00200005fff00000fffd0000ffd100090028001d0016fff0ffee00000000001ffffaffe5ffcf000000000005fff7000000310034ffff00090000, 1024'h0007002100000000ffe800000010000bfff9fff3ffeefff9001b0009fff5fff1001200010008fff1fffa00000004fff90000ffeffff8fffdffef000600230013000efffe000c00130001fffe000ffffb0000ffc0ffdc000f001bffe8ffeffffd000000000018ffeefff9ffec000000000004fffd0000000a0038ffea00080000, 1024'h0000001600000000ffe80000fffc0020ffeb00110020ffee0015ffbbffdbfffa00170027fff0fff8ffe900000013fff50000ffeeffd9ffeefffbfff30019fffb0002fff5fff90001001affe8000400020000ffc4ffec00060017ffd1fff1fff5000000000005fff9000a001200000000000700110000000b002cffda00000000, 1024'h0014001600000000ffef0000001e0014fff80006ffc5000d00350059fff1fff1001dffc90029000300190000001500000000ffec00140005ffe5fff10006ffe8001c00450016000b0006ffd9fff4fff70000ffcfffda0006001b000dffecfff300000000001c000fffdcffa000000000000bfff3000000340032ffecfffd0000, 1024'h0009002200000000ffdc000000130012fff80002ffeefff90023000afffaffec000a0002000afff8fffe0000000800070000ffeb0006fffaffe700050012000700090007000c000bfff20000000400000000ffb5ffce00040027ffe1ffea0002000000000015fff7fffbffed00000000000c000500000005003dffe9fffa0000, 1024'h000c002300000000ffda000000110013fff60001fff0fffa00240008fffcffe9000a00010009fff6fffe0000000700050000ffea0003fff8ffe7000500130007000900070009000dfff1ffff000100030000ffb4ffce00030028ffe0ffe70002000000000013fffbfffbffed00000000000a000700000009003fffe9fffc0000, 1024'h000d002500000000ffda00000015000ffff7fffffff1fffc00240007fffcffe7000a00040008fff6fffd0000000200050000ffea0004fffeffe700040016000900090005000f000effef00030004fffd0000ffb0ffcc00010029ffdfffe70005000000000011fff9fffcffee00000000000c00070000000c0043ffe900010000, 1024'h000c002600000000ffd9000000190013fff60000ffeefffa00270006fff8ffe600100003000afff6fffc0000000600080000ffe800030001ffe6000400150009000a00040012000efff1ffff0008fffa0000ffacffcc0003002bffdeffe70003000000000013fff7fffcffea00000000000d00080000000d0047ffe6fffd0000, 1024'h000d002700000000ffd6000000120017fff40001ffeefff700290008fff7ffe7000c0002000cfff8fffc0000000600040000ffe70004fffcffe200040011000b00070005000c000efff100010008ffff0000ffadffca00020030ffdcffe50003000000000012fff5fff7ffea00000000000f000e0000000a0047ffe6fff50000, 1024'h0010002700000000ffd2000000140016fff30004fff2fffb002a0007fff9ffe5000a00030009fffafffc0000000500040000ffe60003fffcffe10001000c0008000c0009000b000efff40000000200020000ffacffc900040031ffdbffe3000400000000000efffafff7ffea000000000010000a0000000c0047ffe3fff50000, 1024'h000f002700000000ffd0000000180011fff30001fff6fffe00260001fffeffe3000800060005fff9fffb0000000200070000ffe60002fffeffe30000000c0008000c0005000e0010fff40004000300000000ffaaffcb00030030ffdbffe3000900000000000dfffafffdffee00000000001000090000000a0049ffe6fff70000, 1024'h000e002700000000ffd00000001a000efff3fffdfff700000020fffffffcffe4000b00070005fff7fffb0000000200060000ffe600010003ffe4fffe000e0007000b000300130010fff400070008fffa0000ffaaffcd00010031ffddffe3000900000000000efff70000fff2000000000013000b0000000c004affe8fff60000, 1024'h000e002700000000ffd10000001a000cfff3fffbfff50000001efffdfffeffe4000d00060005fff5fffa0000000000050000ffe6fffe0002ffe4fffe000f00080008000000140011fff30007000bfff80000ffaaffd0ffff0031ffddffe3000b000000000011fff90001fff3000000000012000c0000000d0049ffe9fff40000, 1024'h000e002600000000ffd200000012000dfff1fffefff7fffe0021fffdfffaffe2000d00070007fff5fffa0000000300030000ffe6fffdfffdffe50000001100080001ffff000b0012ffef00070008ffff0000ffacffceffff0031ffddffe30009000000000011fff80000fff500000000000f00110000000d0046ffeafff30000, 1024'h000f002600000000ffd3000000100012fff1fffffff9fffb0020fff0fffeffe700080009ffffffeefff80000fffafff80000ffe8fffbfff8ffe5fff8001200080007fffe000d0016fffc00000007fff90000ffaeffd9fffa002fffd9ffe40009000000000008fffdfffdfff200000000000d000d0000000e0047ffecfffc0000, 1024'h000b001f00000000ffd50000000c0022ffef001e0024ffff0000ffb1ffebfff400120013ffd5ffeafff700000007ffe60000ffe7fffa0001fff0ffdf0012ffed0017fff8fff8001f002dfffb000200000000ffbb000dfffd0027ffe2ffe3fffe00000000fff30006000c001100000000000a00160000fffc003cfffc00070000, 1024'h0004000f00000000ffdd0000fff50010ffdd001b006bffeeffcdff78ffe1fff5ffed0029ffaefff2ffca00000005ffff0000fff4ffd1000c0006ffe10010fffcffe7ffc5ffdc0010ffff0019fff0001b0000ffdb003600280016ffedfff6fff800000000ffeeffee001b006800000000000200280000ffde0018000700030000, 1024'h0005000400000000fffc0000ffe6fffcffe3ffc60039fff2fff2ffc5001efffcffd9001bffe5ffecffc80000ffcaffe400000007ffbb00110004000a0009004cffe4ffb3fff6001cffc90010fff80007000000080020001f0002ffe70013fffd00000000fff8fffdfff0002e00000000fffb001c00000013fff7fffa00080000, 1024'h0004ffff0000000000140000ffdb0019ffc9fff500190015006cfffc000d000bfffe0029002ffffaffc90000ffe3ffce0000fffbffd2001afff30018fff60027fff8ffe6ffe50026ffdeffc5ffd0001c00000002ffc20028fff1ffb1001cffe100000000fff9002dffb4ffd400000000ffff002700000043fff8ff8f00060000, 1024'hffeafff800000000001d0000ffcffff8ffc3fff2004000350090ffc40009001800120099003f0014ffad0000ffefffc60000fffdffaa000900070040fff1003d000affc0ffcc001a001affcfffed003800000007ff710041ffd4ff610029fff900000000fff50015ffce000200000000fffe001500000017ffebff30fff70000, 1024'hffcbffdf0000000000370000ffd3ffcffff5fff0002800270070ff9c00190030000d00d6003b001cffb90000ffe3ffdf00000016ffb2ffd900210055ffe600410009ffa8ffe4ffe7005affeb002b00160000002eff630013ffb0ff490036002b00000000ffe6ffea000c003200000000fff3ffdb0000ffcdffc5ff33fff50000, 1024'hffc0ffc600000000004e0000ffe3ffc100440018ffd600060019ffef0015003200080086003a0018000e0000000a00230000002c0036ffd3002a0062ffe2000afff4ffcbfff7ffbb003600280044000100000067ff90ffd3ffa5ffb4002f002e00000000ffe4ffcd0040004600000000ffe8ffc90000ff81ff97ffbcfff50000, 1024'hffdcffba0000000000470000fffdffcb00620022ff9ffff0ffba0048fff800220016fff400200013005a00000034003c0000002f005cffbe002d0017ffebffbdfffa00300012ffa90041001c0038ffe2000000800009ffb2ffb5004b0011001a00000000ffe9ffd70050001100000000ffe1ffad0000ffa7ff9a004f00000000, 1024'hffffffcb00000000002d00000011fff600690023ff91ffb6ff68004bffff000affeeff7cffe1ffdf006b00000019004a0000002e007cffd4001bffda0001ffaeffdb003a0038ffbbffea0025001bffb40000006a008eff8fffe300a7fffd000200000000ffe0ffeb004a000b00000000ffe1ffc80000ffcdffb900dd001e0000, 1024'h002cfff100000000000a00000011004a0022002cffbbffb5ff8b0067ffecffefffe5ff18ffd2ffc6004e0000001300250000000c00780033fff0ffb3000affb3ffd7004900240007ff7efff9ffc0ffce0000003200c9ffc8001e00cafff1ffb200000000ffeb002cffe7ffcc00000000fff600280000003affee00e900270000, 1024'h003a001500000000ffe5000000070048ffc1fff400270013ffef0050ffd9ffe50010ff62ffe5fffc000600000015ffc90000ffe2ffef0061ffe3ffb50008fff100200042ffe50050ffcbffceffaa001e0000fff80083004e002f0079ffefffa2000000000004003fff9bffa000000000000e00470000008500230043000e0000, 1024'h0019001a00000000ffde0000fffbffe9ffb7ffbd004f004300260004fff5ffee00100018ffff0029ffc90000fff7ffbf0000ffe5ff8c001efff8fff0000100360033fffeffd3003b0043fff4fff8003b0000ffe5ffef0078000effeafff7fffe00000000000afff7ffc7ffe000000000000a000900000035002dffa5fff30000, 1024'hfff7000600000000fff80000fff9ffcbfff0ffcf00190012002fffcf0012fffa0001007400160017ffcc0000ffe7fffd00000002ffa7ffd3000b0023ffff003d0008ffcf0002fff00033000c002d00090000ffeeff9d001efff0ff9a0004003300000000fff9ffd90012002100000000fffdffd80000ffec0014ff8ffff10000, 1024'hffedfffe00000000001000000012fff4002b0004ffc4fff10024ffef002100040002003f001fffea00080000ffe8001b0000000d0024ffec00030031000000160002ffdf0034ffdffff20008002bffcb0000fffaffb1ffbffff5ffb90009001e00000000ffeffff60021000900000000fffcffd80000ffdfffffffdd00080000, 1024'hfffd000a0000000000040000001c00210017003effc5fffc00190028fff70005000fffda0011ffe300230000001800110000fff80064001effed00060005ffcf000d001d00150008ffe9fff4fff2ffec0000ffe9ffecffe3000a0009fffaffe80000000000060013fff9ffda00000000000500030000fff1000d000f000a0000, 1024'h000d001a00000000ffec0000000f0015ffef000ffffa000400070028ffe3fff90011ffccfffffff2000500000017fff00000ffed0016001fffebffee0015fff2000d0018fff40027fffafffdffee00130000ffd6000f00280018001ffff2ffe3000000000020ffffffe3ffe100000000000900110000000f0022000bfffd0000, 1024'h0009001e00000000ffe80000000f0002ffecffe300000007000e0013fff0fff5000ffff30003fffcfff300000001ffe80000ffefffdf0009fff2fff8001c001a001200060003001b000bfffb000900040000ffccfff90028001afffffff5fff9000000000025ffefffebffe6000000000009fffb00000019002cffedfffd0000, 1024'hfffe001d00000000ffeb000000130008fff8fff7fff5ffff001bfffefff7fff9000e000d0008fff6fff500000005fffc0000fff1fff1fffffff40009001b00120010fffd000d00090001fff8000cfffa0000ffc3ffda000f0017ffe0fff7fffe000000000023fff4fffcfff3000000000009fff400000005002bffddfffe0000, 1024'hfffb001d00000000ffed0000000c0010fffe0004ffeffff600210003fff8fff900090009000cfff4fffc0000000700030000fff10007fffcfff10013001a000d0006fffd00060006fff2fffd000500010000ffc2ffd200040017ffdffff5fffc000000000023fff5fffdfff7000000000007fffe0000fffc0026ffe5ffff0000, 1024'hfffa001400000000ffec0000fff4001dffed00110019ffee001dffcdffe4ffff000c001efff8fffeffef0000000efff40000fff0ffe2ffe5fffafff90013fffbfffcfffdfff000010016ffe6fffb000d0000ffc8ffe900030012ffd7fff5fff9000000000013ffff00040007000000000006001200000008001fffdffffc0000, 1024'h0009001500000000fff200000024000ffffcfffdffc8000c002c0049fff3fff80020ffd60026fffb00130000001100000000ffee0010000fffeafff70009fff2001c00320020000c0004ffde0000ffeb0000ffcfffde000700170007fff5fff30000000000240005ffe6ffae00000000000effee0000002c002bffebfff90000, 1024'h0001002000000000ffe2000000100015fff90001ffe7fff60025000bfff0fff6001600030012ffecfffe0000000dfffa0000ffec0007fffeffe800070015000900060001000b0012fff7fffa000afffd0000ffb8ffd200080023ffe2fff2fff8000000000022fff0fffaffec00000000000d0005000000060032ffe7fff10000, 1024'h0004002100000000ffe00000000e0012fff8fffdffeafff700230008fff3fff300140005000fffeafffd0000000afff70000ffec0003fffbffe800060019000c0005fffe00090016fff7fffe000affff0000ffb7ffd200080024ffe1fff0fffb00000000001ffff0fffcffef00000000000b0006000000070035ffe9fff50000, 1024'h0004002300000000ffe000000015000ffff8fffdffebfffa00210007fff3fff100150006000effecfffc0000000afffe0000ffec00030001ffea0006001c000b0009ffff00100012fff4ffff000cfff90000ffb3ffd000070024ffe0ffeffffc00000000001ffff1fffdfff000000000000d000200000008003bffe6fffa0000, 1024'h0003002400000000ffe0000000150011fff8fffcffecfff900220005fff3fff000150005000ffff2fffc0000000800020000ffea00000002ffea00080019000c000800000012000cfff5fffe000ffff60000ffb2ffcf00020026ffdeffecffff000000000020fff1fffdffef00000000000f00050000000b003cffe4fff60000, 1024'h0005002400000000ffde0000000d0013fff90000ffebfff100280007fff1ffee000f00060010fff6fffc0000000400000000ffea0003fffaffe600080013000dfffe0000000c000afff10000000dfffc0000ffb1ffccffff0029ffdeffec000200000000001dffeffffbffef00000000000f000d0000000a0038ffe8fff10000, 1024'h0007002300000000ffda000000130011fff8fffeffeafff900280008fff5ffed001200080010fff1fffe00000006fffd0000ffea0004fffdffe600040010000a0006000200100010fff4fffe000bfffa0000ffb1ffcb0001002affdeffed0001000000000019fff3fffdffeb00000000001000080000000c003bffe7fff10000, 1024'h0007002400000000ffd80000001b000ffff8fffcffe9fffd00230005fff8ffed00170008000effeafffd0000000800000000ffe900050003ffe6000300130009000bfffe00160015fff50001000efff50000ffaeffcc0004002affdcffec0001000000000019fff10001ffee0000000000100003000000090041ffe6fff20000, 1024'h0007002700000000ffd80000001b000ffff7fffbffebfffd001f0001fff5ffee001a0007000bffe8fffc00000008fffd0000ffe800020004ffe7000100190008000bfffd00160016fff600010011fff30000ffaaffd00004002bffddffeb000000000000001dfff00001fff000000000001000050000000a0044ffe8fff40000, 1024'h0007002800000000ffd9000000150010fff4fffcfff1fffa001ffffbfff4ffee001600080009ffeafff800000006fffd0000ffe8fffd0001ffe80002001a00090004fffa00110014fff30001000ffff70000ffaaffd10004002bffdbffea000100000000001ffff10000fff500000000000f000c0000000a0043ffe7fff30000, 1024'h0007002700000000ffdb0000000c0010fff3fffdfff6fff80022fff8fff6ffee0011000b0008fff1fff700000002fffa0000ffe9fffafffaffe800030018000c0000fff9000a0013fff40001000dfffd0000ffaeffd10001002affd9ffea000400000000001cfff6fffdfff600000000000e00130000000a003fffe7fff30000, 1024'h0008002400000000ffdc00000008000bfff30002fff9fffe0021fffefffbffec0009000a0008fffafffa00000004ffff0000ffea0000fff6ffe90006001300070001ffff0002000ffff50006000700070000ffb7ffcd00010027ffdcffe70008000000000016fffbfffcfff800000000000c001300000002003bffe7fff40000, 1024'h000c002000000000ffdd00000004000efff000080006fffb001dffe7fffeffed0001000dfffafff9fff50000fff9fffa0000ffecfff5ffefffecfff8000f0001000100000001000d0002fffdffff00030000ffbcffdefff90023ffd9ffe6000c0000000000070006fffdfffb00000000000900100000000a0038ffe9fffe0000, 1024'hfffe000d00000000ffe10000ffe6001effc800180070fff10016ff5fffe4fff2fffd005fffd1fff9ffb600000007fffd0000ffefff9dffec000bfff0000d0000ffe3ffc8ffe3fffdfff4ffddffdc00180000ffc5ffee00180010ffa6fffdfff300000000fff100130015004f000000000003002900000014001effb7ffff0000, 1024'hffdefff40000000000090000ffc6fff0ffcfffc2007ffff30029ff4700230002ffde00bffff5fff6ff890000ffd5fff90000000eff6afff10026004b00070072ffc8ff5dffe6fff5ffb00001fffa001c00000005ffb20025ffe2ff610031000500000000fff0fffb001f008a00000000fff600230000fffcffddff7efff60000, 1024'hffc9ffd40000000000440000ffc2ffdbfff4ffc7001800200080ffc0002c0026001300cb005d0018ffc20000ffeaffe40000001bffa0ffda00280076ffec005ffffaffa0ffecffe20009ffd8001a001600000044ff510005ffadff4f0043001000000000fff200070006001f00000000ffeffff100000001ffafff39fff00000, 1024'hffbcffc100000000005d0000ffd5ffc400360014ffc800180060fff00020003e001500ae0062001e00040000fffe00070000002c001affb90028006affdb000f0002ffd9fff9ffba0059fff7003ffffd00000066ff55ffc6ff96ff790037003400000000ffdfffea0028001800000000ffe7ffbd0000ffa5ff98ff70fff90000, 1024'hffccffb80000000000550000fff8ffd3006c004dffa6ffefffd4001a0003003400090021001f0010005100000021003f000000330087ffcc002a002cffdcffb8fff70014000dffa4004a0027003dffde00000082ffecff96ffa900180019002800000000ffd3ffdd0052002b00000000ffe5ffb90000ff7cff8e003000060000, 1024'hfffcffc800000000003400000012fff3006a0044ff9bffc9ff610060fff50014ffe8ff66ffdbfff400740000001e00490000002c00a6fff40017ffd6ffecff96ffe3004b0021ffc1fffb00330010ffc90000007c00a1ff9fffdd00c3fffeffff00000000ffdfffed0038000900000000ffe7ffd40000ffb3ffa600e700180000, 1024'h002effea00000000000700000015002e00210026ffd5ffd5ff580061ffe9fffaffe8ff05ffafffd3005a0000001600080000000d0066002bfffdff8b0006ff99fff4006300120016ffcefffeffc4ffda0000004a0108ffdd001200faffecffbf00000000ffed002dfff1ffcd00000000fff200110000002effe0010a00290000, 1024'h003d000d00000000ffea000000050036ffcefff70035fffbffa10038ffe2ffe7ffecff40ffb5ffe2000500000005ffd70000fff1ffff0060ffeeff9f0016ffe6fffd002cffe40053ffb4fff6ffa700180000001000d20049002600adfff0ffab00000000ffff0030ffb5ffd50000000000000047000000620010009300210000, 1024'h0029001600000000ffeb0000fff60004ffadffac004c002e0018002effecffe7000affd500010022ffcb0000fff4ffbe0000ffe8ff8b0044fff4ffe6000a0042001b0006ffd70044fff9ffe9ffdd00360000fff600260080001400210000ffd90000000000120007ffa6ffc700000000000a002b0000006d0022ffd3fffe0000, 1024'h0000000a00000000fffc0000fffdffd1ffeaffb3fffd00350053001d0011fffe00180053003a0035ffe20000ffe5ffd60000fff9ffa9ffeafffc0023fff2004c0033fffbfffd0005005efff70036000f0000fff7ff93002ffff8ffaf0003002c000000000003ffe0ffe2ffcf000000000007ffd900000013001aff7dffec0000, 1024'hfff2fffb0000000000000000fffafff300080026ffebfff3003fffc9000f0004fff700610019fffcffe60000fff5002200000005ffffffc3fffd001affeefff6ffefffe90010ffd70016fff3000efff10000ffe9ff92ffddfff5ff900001002700000000ffe3fff6001a001a00000000fffaffdc0000ffd4000bffa4fffa0000, 1024'hffeffff40000000000060000ffe30026ffec001e0039ffe10028ff7a00130003ffe90064fff4ffd8ffca0000fff7001000000007ffe0fff5000e0021fffe000effd5ffb0fffdfff0ffadffe3ffd500000000fff8ffd2ffe4fff4ff950017ffec00000000ffde0029001a004e00000000fff9002100000002ffeeffc100070000, 1024'hffebfffc0000000000220000fffefff60008ffe8fff60025003c001500300014fffb0032002c0006fff80000ffe0ffe900000009001e003500000049fff6003c001affd4ffff0015ffe3000e000900080000001dffbd0003ffe4ffca002000020000000000010013ffe4fff3000000000004000b0000fff3ffe0ffc100080000, 1024'hffff00080000000000190000001affe80003001dffab0039005e0091000100150013ffdd0051001f00170000fffffff60000fff8004a001effe20012ffecffe50029004c0002000f0035ffebfffe000a0000fff9ffa8001dffeffffa0004000b0000000000230001ffb8ff8c000000000009ffd90000fffe0006ffb200000000, 1024'hfffe001500000000fff7000000110000fff5000fffdf000e0038002bfff50003000ffffb0023ffff000000000009fffc0000fff2000cfffbffee00010009fff1000b0022000600090011ffe9fffa00040000ffccffc7000e0009ffe7fff9000300000000002a0000ffe9ffcf00000000000affef0000000b0020ffcefff80000, 1024'hfff4001900000000fff10000000e0009fffefffdfff8fffa001cfff0fffaffff000e001a000afff4fff70000000300000000fff4fffafffefff800110018000f0003fff3000e0003fff5fffb000dfff70000ffc4ffd5fffe0012ffd8fffd0001000000000027fff70007000100000000000bffff0000ffff001fffe1fffa0000, 1024'hfff3001700000000fff30000000d000dfffd0004fff6fffa001dfff6fff70003000b0014000bfff6fff70000000700010000fff4fffffffffff60010001400090001fff9000a0001fff5fff70007fffb0000ffc7ffd700030012ffdcfffffffd00000000002bfff70002fffe00000000000bffff0000fffb001affe0fff70000, 1024'hfff4001700000000fff300000007000bfffdfffefff1fff900200003fffc00030008000d0010fff4fffa00000003fffc0000fff50002fffcfff300120015000ffffefff900050009fff0fffa000400010000ffc9ffd600040012ffe00000fffd00000000002ffff8fffdfff800000000000a00020000fffe0017ffe5fff70000, 1024'hfff4000f00000000fff30000ffee0019fff0000c000bfff10022ffe0ffed0007000d00180006fffbfff50000000bffef0000fff3ffeeffe3fff70000000ffffefff6fffdffec00080013ffe9fffd00100000ffd1ffe5ffff000dffd9fffbfffb00000000001cfffefffeffff0000000000050014000000030014ffe2fff60000, 1024'hfffe001500000000fff60000002b0003fffffff7ffcf0012001e003afffbfffe001effdf0020fffb000e0000000d00080000fff0000b0016fff2fffe000cfff5001b0025002700070001ffe50008ffe40000ffcfffe2000600110004fffafffa0000000000330004fff2ffbf000000000010ffe9000000200024ffeafff60000, 1024'hfff8002000000000ffea0000000b000dfffbfffeffe7fff80021000bffeffffe001700030015ffecffff00000008fff40000ffee0004fffdffed0009001b0009fffe0000000b0010fff5fff9000dfff90000ffb9ffd60001001effe5fff7fffa000000000035fff2fffbffef00000000000f0006000000090026ffeaffee0000, 1024'hfff9002200000000ffe800000011000afffcfffbffe7fff900210007fff1fffb001800080012ffe6fffd00000007fff40000ffee00040000ffee000a0020000c0001fffa000f0015fff4fffc000ffff70000ffb4ffd40005001dffe3fff8fffb000000000033ffef0000fff100000000000d000200000007002bffeafff40000, 1024'hfff9002300000000ffe800000013000ffff9fffcffe8fffa00200005fff0fffd001900070012ffe8fffc0000000efff70000ffed00020000ffee000a002200090005fffd000f0012fff7fff90010fff80000ffb3ffd30007001effe1fff6fff9000000000035fff1fffffff000000000000e0004000000040031ffe5fff30000, 1024'hfffc002300000000ffe80000000c0010fffafffdffecfff500210002fff0fffc001400080010ffedfffa00000004fff70000ffed0000ffffffeb000a001f000dfffefffb000c000efff4fffd000ffff80000ffb3ffd200010021ffddfff4fffd000000000030ffeffffcfff500000000000f000900000008002effe5fff50000, 1024'hfffb002200000000ffe70000000c000ffff9fffeffedfff400280004ffeffff80014000a0013fff2fffa00000002fffa0000ffed00020000ffeb000a0019000efffafffb000c000efff1fffc000efff90000ffb1ffd000000021ffdefff6ffff00000000002dffeffffbfff1000000000010000d0000000b002effe6fff40000, 1024'hfffb002300000000ffe400000015000bfffbfff8ffe4fffe0025000bfff2fff9001c000a0016ffeafffe00000006fff40000ffec00060005ffea0009001a000e0007fffc00140016fff9fffd0015fff20000ffb2ffce00040023ffdffff6fffd00000000002cffecfffcffeb0000000000110003000000080033ffe5fff10000, 1024'hfffd002600000000ffe10000001b000cfff9fffcffe2fffe00220009fff0fff9001f00060014ffe1fffc0000000cfff70000ffea00060007ffe90006001f00080009fffc00170019fff8fffc0013fff10000ffacffce00090024ffdefff3fffa000000000031ffedffffffed000000000011ffff000000070039ffe2ffef0000, 1024'hfffc002900000000ffe1000000150011fff6fffbffeafff90023ffffffeffff8001c00090010ffe4fff80000000bfff50000ffe9fffd0002ffea00090025000e0005fff800110017fff3fffa0011fff60000ffa7ffd000080026ffdafff2fff9000000000036fff1fffefff2000000000010000600000009003affe1fff10000, 1024'hfffb002800000000ffe20000000b0011fff60000fff1fff80024fffdffeefff80015000b000efff0fffa0000000afff60000ffe9fffefffaffeb000b0022000c0002fffc00050011fffafffd000f00000000ffabffce00040025ffdaffeffffe000000000033fff1fffdfff500000000000f000c000000030036ffe2fff20000, 1024'hfffe002400000000ffe200000002000efff60004fff7fff20021fffcfff2fff50006000a000afff9fff900000004fffd0000ffecffffffefffeb0009001a0009fff8ffffffff0008fff70002000800070000ffb3ffd0ffff0023ffddffec0005000000000028fff3fffdfffc00000000000d00100000ffff0031ffe8fff40000, 1024'h0005001f00000000ffe30000fff70015ffe900050007ffed002cffeafffefff0fff600110006fff8ffe90000fff800000000ffeeffeeffebffeb00070012000cffe9fff6fffb0006ffdcfff6fff2000c0000ffb8ffd0fffd0021ffcffff000030000000000190008fff50000000000000009001d00000010002dffdefff90000, 1024'h0004001900000000ffea0000ffe3001dffceffff002dfff90052ffc1000bfff2ffee003e000cfff7ffc70000ffe8fff00000ffefffc8fff4fff00014000a0021ffe3ffd9ffed000fffc8ffdfffd900190000ffbfffb600090017ff9dfffffffa0000000000080022ffe400090000000000070030000000290024ffa7ffff0000, 1024'hffe6fffe00000000fffe0000ffcc0012ffbb00020088001c005eff43fffa000c001000bcfff80010ffa00000fffaffd00000fff4ff74ffe70018001d000000280002ffadffc900060029ffc3ffe500300000ffe0ffa40024ffeaff530018fffc00000000ffea002500060046000000000000002400000018ffffff4effff0000, 1024'hffb8ffd400000000002e0000ffc9ffbd0004ffed00760014000cff3400170029fff600fefff20020ffaf0000ffeeffff00000021ff9effd40044005cfff2004afff0ff6affcfffd000460028003a002400000042ffa1000fffabff5e0038003600000000ffd9ffcd005600b100000000ffebffe90000ff89ffaaff75fff80000, 1024'hffc0ffb100000000005d0000ffe7ffac0069fffdffc5fff4ffbffffb0022003afff900520017001800310000fffb002700000041003cffbf003e0046ffe10006fff6ffd90009ffa90055003f0060ffe20000009ffff3ffb3ff960005002f003f00000000ffd8ffbd005d004f00000000ffdbffa90000ff72ff76002200030000, 1024'hfff2ffb400000000004f0000000bffe80083004dff71ffceff6e0088fff50025fff8ff6cfffcfffd00900000002e004b0000003800c5ffde001dffe6ffe3ff86ffeb00610021ffaf001d00300022ffc7000000a20084ff8affc300c50005000600000000ffd8ffe6003ffff500000000ffdfffbf0000ffa0ff8b00e000160000, 1024'h002cffd80000000000160000001c00270041003bffb0ffbfff420084ffe2fffcffe4feefffb9ffe100760000002300340000001a0090001e0001ff8dfff5ff80ffe3007a0022ffecffc7000fffd2ffca00000066010bffbd00080118ffebffcb00000000ffe2001a0005ffd100000000fff0000000000015ffcc012d00230000, 1024'h0042000100000000ffe90000000b003effdcfff60020ffecff86004cffe9ffe1ffe3ff1bffb1ffe6001b00000007fff10000fff700090056fff0ff8f0006ffd3fff30045fffc0039ff99ffebff9fffff0000002000f00028002f00d1ffeeffa800000000fff8003effbeffc8000000000002004200000074000600c1001d0000, 1024'h0032001700000000ffe20000fffb000fffb0ffb5004a00390000002d0004ffe60003ffb2ffea000dffdf0000fff0ffb00000ffe6ffa40046ffefffd1000b002c002b0014ffd7005dfff5ffe5ffc600340000fffa0050006e001c003bfff7ffd2000000000008002effa5ffbc0000000000060030000000720025ffff000c0000, 1024'h000c001000000000fff40000fffeffd6ffd0ffcb00300040003d0004fffefff4001400410018002effd10000fff5ffd70000fff1ffa100060001000d00030034002dfffaffe1001b004dfffc0010002c0000ffedffb80055fff8ffc5fffc0018000000000002ffecffddffe9000000000002ffed000000180024ff88fffe0000, 1024'hffebfffa0000000000060000fffcffdd0001ffe9000cfff50032ffb50003fffe0004008300170010ffce0000ffed001b00000009ffb5ffcf00130028fffd002efff4ffc90018ffce0020fffb002fffea0000fff0ff97fffdffebff8d000e002b00000000ffeeffd20026002e00000000fffbffd10000ffea0007ff91fffa0000, 1024'hffe6fff30000000000160000fff2000f00220000ffceffd40030ffd80027000dfff3004b0025ffd9fff90000ffe30014000000120021ffe6ffff003dfff70024ffe0ffbf0028ffe4ffc6fffe001affd400000009ffb1ffb9fff3ffa80019000a00000000ffe5fffc001b001900000000fffa00000000ffe5ffe9ffdffffe0000, 1024'hfffbfff00000000000110000ffec002bfff5003bfffd000a003ffffaffe900100024001c0021fff100040000002cffee0000fffb0024000bfff9000ffff1ffd900050007ffe1000effffffd6ffdc001d0000000effd00002fff1ffd9000cffd500000000ffeb0024fff0fff100000000fffd001f00000007ffebffcafff80000, 1024'hffe9ffe400000000000f0000ffeaffe2ffe6ffee005500120005ff96ffed000f0011007cfff6000fffc40000000efff90000000cff99fff10027000ffffa001cfffaffc2ffe4ffef002cfff8000b00180000001dffe00033ffd7ffb80021000500000000ffefffe20024005100000000fff7ffeb0000ffeeffddffa5fff50000, 1024'hffd5ffdf00000000003300000001ffca0031ffb2ffc8ffeb000800030042001bffe800570034ffefffed0000ffcc00210000002bfff7fff4001a005afff70060ffe6ffa7003cffd3ffc900240043ffc80000003effb8ffe0ffceffbf00380024000000000001ffca0024002b00000000fff4ffc50000ffd0ffc1ffdafffc0000, 1024'hffeeffee000000000034000000190016002c001aff69000e005d009b000800200037ffd60074ffec00410000001f000700000008006e0013ffed0030fff4ffe1001c00420030fff6ffe7ffc80002ffd700000018ffa3ffd1ffe7fffc0019ffde000000000021001dffdaff83000000000003ffdc0000001dffe1ffdafffa0000, 1024'hfff4000b000000000008000000140015fffe002bffc5000d0047003dffe600140027fff20037fff3001000000022fffd0000fff4002e0007ffed00050006ffd8000e003000090008000dffd3fff4fffc0000ffd6ffc000040001ffe90005ffeb0000000000320008ffe4ffbc00000000000bfff00000000b0010ffcafff30000, 1024'hffeb001600000000fff70000000a000cfffefffcfff6fff7001bfff4fff5000d00100019000effeffff400000006fff80000fff7fffb0000fff80013001700140002ffef00090008fffbfff8000efffa0000ffcaffdb000a000dffd90007fff9000000000035ffed0001000200000000000cfffb0000fff60013ffdefff20000, 1024'hffea001400000000fff900000008000dfffe0000fff4fff7001dfff9ffef000e001500150011fff1fff70000000afff70000fff6fffc0000fff800100016000d0000fff500080007fffcfff2000bfffa0000ffcbffdc0009000cffde0008fff5000000000038fff00000fffd00000000000dfffd0000fffd000effdffff00000, 1024'hffe9001400000000fffa0000000600080000fffaffedfff6001d0001fff5000e001200130016ffeefff900000007fff60000fff80000fffcfff8001500160012fffcfff200070009fff7fff8000ffffc0000ffceffda0007000affe00009fff900000000003bffed0000fffc00000000000bfffd0000fff8000cffe4ffed0000, 1024'hffef000d00000000fffb0000ffe70017fff80009fff6ffea0021fff3ffed000f000f000e0012fff1fffc0000000cffe90000fff7fffbffdefff6000800100001ffedfffaffeb000b000effec0005000f0000ffdcffe5fffc0009ffe10000fff8000000000028fff6fffcfffa00000000000200150000fffb0007ffecffeb0000, 1024'hfff7001500000000fffb00000028fffcfffdfff6ffe1001c00180028000a00040011ffe900170002000700000003000a0000fff10005001afff80007000cfff8001b001c00210003fffdffea0002ffea0000ffd3ffe30004000afffbfffc000200000000003b0010fff5ffcf000000000010ffec00000017001affe3fff90000, 1024'hfff2002000000000fff4000000050002fff90005fff300010024000bfff70005000700040012fffefffc0000fffcfff50000fff10004fffcfff2000c00190005fff9000700010008fff5fff9000300030000ffbcffd7fffe0014ffe6fffb00050000000000430001fff4fff00000000000100009000000050019ffe5fff40000, 1024'hffef002200000000fff100000015fffefffc0000fff10009001f0009fffb0002000c0007000ffff9fffd00000000fffc0000fff000050006fff6000f001d000700060004000d000afff5fffa0007fffa0000ffb7ffd600030014ffe6fffc0004000000000045fffefffcfff0000000000010fffb000000010020ffe4fff80000, 1024'hffef002300000000ffef000000110008fffc0000ffedfffd001f0007fff40004000f0004000ffff3fffd00000008fffa0000ffee0003fffdfff3000e0022000600020003000a000bfff9fff70009fffd0000ffb3ffd700060016ffe6fffaffff000000000048fff6fffffff000000000000effff0000ffff0023ffe7fff40000, 1024'hfff1002300000000ffee00000009000dfffd0000ffeefff0001f0001ffea000300130009000fffeefffb00000008fff60000fff00000fff9fff2000d0025000cfff9fffb0007000bfff3fff9000dfffd0000ffb1ffd800040019ffe4fffcfffa000000000044ffee0000fff800000000000e0006000000020022ffebfff40000, 1024'hffef002100000000ffee00000012000dfffffff9ffeafff4001e0002ffeb0003001b000c0013ffedfffc00000009fff90000fff0ffff0002fff3000e002100100000fff90013000afff5fff80015fff10000ffb3ffd70003001affe2fffefff9000000000040ffe90002fff50000000000110000000000050025ffe8fff10000, 1024'hffef002400000000ffec00000015000cfffffffbffe0fff7001f000afff10005001900060016ffe9fffd0000000afffa0000ffef00060001ffef000f0020000d0003fffb0016000dfff2fff70015fff00000ffb1ffd30004001dffe1fffdfff9000000000046ffeefffeffef000000000012fffe0000ffff0028ffe6ffeb0000, 1024'hfff2002700000000ffe90000000f000dfff80001ffea000000220009fff30004001700030014ffebfffe0000000dfff40000ffeb0004fffeffee000d0023000500060003000a0012fff4fff50008fffd0000ffaeffd00005001effdffff6fff8000000000049fffcfffaffef000000000012000400000004002affe1ffec0000, 1024'hfff2002800000000ffea000000090006fff70003fff7fffd00210000fff7000000080008000dfffcfffa00000004fffc0000ffecfffefff5fff1000f00210007fffd000300020007fff6fffd000700060000ffadffd00000001bffdefff20007000000000048fffefffdfff8000000000011000a0000fffe0029ffe2fff00000, 1024'hfff6002500000000ffeb0000fffc000cfff100070000fff2002afff3fffbfffcfff7000d0009fffeffef0000fff5fffe0000ffeefff6ffeeffef000d001b000affeafffdfffe0001ffe3fff6fff900070000ffaeffd0fff9001dffd5fff5000800000000003c0005fff6fffc00000000000e0015000000080024ffe0fff70000, 1024'hfff8002000000000ffed0000ffe7001affd80005001dfff3004affd50005fffcffee0029000efff8ffd40000ffecfff20000ffeeffdcfff0ffef001400130017ffdeffe6ffee000dffcaffe2ffde00180000ffb2ffbf00040017ffb10000fffc00000000002c001cffe6000100000000000b002e0000001d001fffbcfff90000, 1024'hfff1001400000000fffb0000ffcd0015ffc3fff8003f00070078ffb3000c0003fff6006e00220001ffb40000ffe6ffda0000fff1ffb3fff0fff7003000090036ffe1ffc3ffd50016ffd7ffd6ffda00310000ffc7ff8e001c0001ff740011fffa0000000000160021ffdb0010000000000005003800000023000eff71fff70000, 1024'hffddfffc0000000000160000ffcaffecffdcffef003700210082ffb000140013000800b20039001fffbc0000ffedffdc00000000ffb2ffdd000c0052fff90042fffaffb7ffcffffe001dffea000800360000fff6ff5c0019ffd9ff55001f001a00000000ffff0004fff7002100000000fffc00120000fff2ffeeff46fff30000, 1024'hffcbffd900000000002f0000ffe1ffd100220014000f0017002dff9e0007002c001900b000190021fff500000000fff500000019ffebffba00280038ffea00090014ffd2ffe9ffce008b00030043000600000034ff98ffddffb9ff88001d003a00000000ffd8ffdd003e003f00000000ffeeffca0000ffa3ffc6ff9100000000, 1024'hffd1ffc200000000003700000003ffd6006d004affe0ffd9ff7cffc1fffa002dfff60021ffcafffb004000000018003c000000320073ffd200310006ffecffbdfff3ffeb0009ffb4005a004e004affd8000000710049ffa7ffbe00360011002d00000000ffc3ffbd0078007600000000ffe2ffbe0000ff52ff9f007600130000, 1024'h000effcd00000000002600000017000c00630038ffacffaeff270059ffee000fffdaff2affb0ffcf006e00000017003e0000002c00ab0018000effb6fff9ffa0ffd500370021ffe5ffd200450001ffc40000007e00fdffb8fff100fcffffffe100000000ffdaffe1002f001a00000000ffe5ffec0000ffbcffac013200220000, 1024'h0046fff500000000fffd00000013004dfffe0006ffd6ffd3ff740099ffd6fff0fff7fed4ffc3ffc9004900000018ffe900000001004f0059ffe6ff80000affb9fff4006800090043ffa3ffeaffabffea0000003d0119001800270112fff3ff9200000000fff9002affb5ff9b00000000fff900310000006ffff3010300230000, 1024'h0042001600000000ffde00000000003bffa8ffc90039001afff00049ffd6ffe80016ff6fffe6ffefffe800000009ffa80000ffe2ffb90062ffe1ffa8000e0011001e002bffdd006fffe3ffceffb500260000fff8008b007d002e0070fff8ffa20000000000070023ff8effa000000000000b004400000094002d002c00080000, 1024'h0015001400000000ffe60000fff7ffeaffbbffa8004500420033fffefff3fff60029003800110020ffc40000fffaffaf0000ffe9ff7e001cfff8ffff0006004f003affe8ffd800410051fff5001300330000ffedffd8007b0008ffcf0001fffb000000000001ffe4ffcaffe4000000000008000500000034002cff8cfff00000, 1024'hfff7000000000000000100000003ffc4000effd9ffe50016002bfffb00140000000f006500270014ffed0000fff0000000000007ffdbffcd0004002cfffc00310017ffe10008ffee0054001e004affff0000ffffff91000cffedffa9ffff003e00000000ffefffc20018000e00000000fff6ffc20000ffc90012ffa1fff50000, 1024'hfff8fff4000000000007000000100001002f002affcbffe0fffaffeb0000fffe0006001e0005fff1001c0000001000340000000c0031ffd30006000b0000ffdefffa00050027ffcb000a0007001effd400000001ffd8ffb9fffbffe4fff6001600000000ffdefff00036001700000000fff7ffd70000ffd200050009000b0000, 1024'hfff6fff000000000fffb0000000b0020000d002b002bffdbffc3ffa1ffe1fff900070011ffccfff3000100000027003500000004fffc0003001affee0003ffd7fff0ffee0012ffd3ffdffff8fff3ffe5000000030031ffdf0003000affffffe600000000ffe50007003e004b00000000000100050000fff6fff5002a00060000, 1024'hfff0ffef0000000000060000fff6fff00008ffcd0020ffe7ffccffd9000cfff9fff20019ffeefff9ffec0000fffa00190000000fffd30006001b001c00030032ffe0ffc0000affedffbc001b000cfff800000021001d0009fff5000b0017fff8000000000002ffe60026004500000000fff900030000fffaffd90020fff40000, 1024'hfff3ffe90000000000190000fff4fffe0009ffd9ffe0fffc0019000bfffe00100026001b0026ffed000600000006ffdf0000000dffd9ffe50010000a000000180009fff9001000010019ffd60015ffea00000023fff3fff9ffe5fff2001bfff1000000000001fffd0006ffe000000000fff5ffe300000026ffdfffeafff60000, 1024'hffdbffe200000000001b0000000700050020001e0007fffaffdeffa8ffd9002700380049ffefffde00090000002bfff0000000100005fff90022fffd0007ffe7001affde000afff50055fff4002effdf000000260014fff1ffdbffea001bffee00000000ffe9ffdf003f003700000000fff8ffd90000ffccffd8fffafffe0000, 1024'hffdcffe20000000000210000000cffe90026fffbfffaffd0ffa3ffe0ffee001bfff9000cffecffd5fff1000000130036000000200014001d0020001a000b0010ffd1ffb5001fffdfffbf00320023ffdb000000380032000fffdf0020002affea000000000010ffb70039006900000000fff8ffe20000ffb5ffbf0034ffef0000, 1024'hffeffff100000000002b0000000d0000001cffb3ff9efffb0004007b000f001b0025ffbe0047ffe0002400000001ffe700000011000300180005001e0010002e000d001000360007ffcaffdc0016ffcd0000002d000efff8ffed00340026ffd50000000000430005ffe4ffad000000000002ffde00000044ffcf001affee0000, 1024'hffea000600000000001900000012001300060014ffb00013004a005affe300210038ffe6004bfff4001d00000022ffe60000fff70027000dfff2000c000bffe5001a00390012000a0018ffc30001ffef0000ffe8ffc80000fff8fff90010ffe0000000000048000cffdbffa000000000000effe800000023fffaffccffec0000, 1024'hffe000130000000000010000000b00080003000bffe7fff400240000ffe8001a00150019001bffecfff60000000cfff80000fff9000a0001fff8001500150008fffafff5000900030002fff30011fff80000ffcaffd3000b0004ffda0010fff7000000000048ffe40000fffd00000000000ffff30000ffed0004ffd6ffe80000, 1024'hffde001200000000ffff00000008000e0002fffaffeefff40019fff7ffec001a001c00170016ffe8fff90000000dffef0000fff9fffa0000fffd001400190011fffffff0000b0007fffdffec0012fff40000ffcdffe300070007ffe00012ffef00000000004cffec0004fffe00000000000ffff80000fffb0001ffe2ffe70000, 1024'hffde001200000000000100000006000b0005fffeffe7fff300190002ffee001b001800110019ffe7fffc0000000dfff00000fffa0006fffefffa001700190010fffafff10007000afffbfff40012fff90000ffd0ffe100080006ffe40011fff200000000004effe80002fffe00000000000dfff90000fff1ffffffe7ffe50000, 1024'hffe8000c0000000000000000ffdd0019fffc0009ffeaffdf001f0005ffea0017000cffff0019ffee00020000000fffe60000fff90007ffd7fff3000c00130002ffe0fffbffe2000f0007ffef000500170000ffdfffebfffd0007ffee0005fff400000000003bffeffff8fff6000000000001001c0000fff3fffbfffbffe30000, 1024'hfff2000f00000000000300000019fff00000ffeffff100240015001900210008fffffffc0012000e00040000fff300090000fff7ffff0011ffff0017000800040018000f0013fffdfffbfff6fffffff70000ffe4ffdcfffaffffffeeffff0011000000000036001bfffaffe200000000000bfff00000000a0008ffde00000000, 1024'hfff000170000000000010000fffffff7fffa0015fffa000a0028001400020008fff1000200130018ffff0000fff500050000fff7000ffff5fff7000e000dfff5fff2001afff8fff4fff6fffafff3000e0000ffccffd2fff30006ffeafffb001400000000003e0012ffefffef00000000000e00080000fffd000bffe1ffff0000, 1024'hffed001a00000000fffa00000018fff6fffd0002ffff001400190004000e0004fff500080007000ffffb0000fff2000c0000fff50001000bfffd0011001100020005000d0011fff5ffe9fff8fff8fff80000ffc4ffdbfff7000cffe8000000100000000000430014fffcfff4000000000012fff7000000040011ffe200020000, 1024'hffe8001e00000000fff700000016fffffffd0002fff6000c002200070004000800030006000d0001fffd0000fffb00020000fff100050008fff900130019000400050008000b0004fff2fff3fffcfffd0000ffb8ffd80000000dffe6000200070000000000500008fffdffed000000000010fff9000000020014ffe2fffd0000, 1024'hffe5002100000000fff50000000f0009fffc0003fff2fffc00230004ffef000d000f000a0011fff6fffb00000007fff60000fff100040000fff6001000220009ffff00020006000afffafff30007ffff0000ffb1ffda00080011ffe50004fffc000000000055fff4fffcfff2000000000011fffe0000fffc0019ffe4fff50000, 1024'hffe4002200000000fff300000015000dfffffffdffecfff6001b0000ffea00100017000a0011ffedfff900000009fff70000fff100000007fff5000f0023000f0002fffa00120009fff8fff30012fff10000ffb0ffde00090016ffe30006fff6000000000057ffeafffffff6000000000015fff90000fffd001bffe4ffed0000, 1024'hffe4002200000000fff10000000b0011fffcfffeffebfff6001e0008fff00011001100040015fff2fffc0000000efff60000ffef0003fffcfff10014001f000cfffeffff00060009fff4fff3000b00000000ffb3ffd900090018ffe40002fff600000000005cfff2fffbfff400000000001400040000fff80018ffe5ffe40000, 1024'hffec002200000000fff00000fffa000ffff20006fff7fff700280003fffa000effff00050012fffafff600000003fff30000fff0fffaffe9ffef000f001b0007fff30006fff50007ffefffeffff800110000ffb4ffd400030017ffdbfffdffff0000000000560006fff1fff4000000000010000d0000fffe0017ffdeffe90000, 1024'hffef001f00000000fff30000ffe60016ffdc000b001cfff50041ffde000a0008ffe2001e000d0002ffd90000ffebfff90000fff1ffe2ffe9fff1001500120010ffdcfff4ffea0001ffcdffe3ffd8001c0000ffb4ffc5ffff0013ffb8000100020000000000430020ffe4000300000000000e0025000000110014ffc0fff60000, 1024'hffe8001800000000ffff0000ffd20010ffc8fffe0041000a006effbd00170009ffe3005b001b0010ffbb0000ffdcffe70000fff2ffbefff3fff90030000a002effdeffd3ffd90009ffc7ffd6ffcd002f0000ffbfff9a000f0001ff83001200010000000000320033ffd8000d00000000000c0036000000220005ff80fffc0000, 1024'hffd700050000000000160000ffcaffefffd3fff5003c0027008bffbd001e0016fff6009b00390027ffbb0000ffe2ffde0000fffbffb8ffe400080052fffb003cfff2ffc6ffca00000006ffe0ffef003e0000ffe4ff620017ffddff5d001f001a000000000020001cffe60012000000000002001c0000fffeffecff49fff50000, 1024'hffcaffe900000000002d0000ffceffcc00070006000e001b0063ffcd00130022000200a9003f002fffe10000fff5fffb00000011ffe2ffbd001b0057fff00021fff4ffd2ffd7ffd50044ffff0023002800000018ff5ffff3ffc0ff7400200037000000000004ffec0018002900000000fff4ffe90000ffbdffccff6afff40000, 1024'hffd1ffd30000000000380000ffedffce00510021ffc0ffeefff9ffff001000210000004a00210015002f000000070029000000260048ffb300200038ffedffedfff2fff80005ffb6004500270043ffef0000004bffc2ffacffc0ffe50011003a00000000ffe4ffd40049002d00000000ffe8ffc50000ff90ffb7000500030000, 1024'hfff9ffd60000000000260000000e0007005c0050ffa7ffc4ff930027fff10013fff4ffa1ffe0ffe6005d000000180039000000220092ffe5000effdbfff3ffa0ffe800340023ffca000e001e0015ffc400000050006eff96ffe90079fffb000300000000ffd4fff1003a000d00000000ffecffdc0000ffb8ffc600ac001a0000, 1024'h0024fff200000000ffff00000017003f001b003affecffc8ff70002affdefffbffecff3affabffc5003d00000015000e00000008006b0041fff7ffa00004ffacffec00330010001bffbc0009ffcaffdb0000003000e7ffe8001900c3fff4ffb800000000ffe10019fff7fff600000000fff9002000000014ffea00e200220000, 1024'h0035001100000000ffe700000011002fffd0ffe000240008ffb8004effdaffeb0008ff54ffcfffde00030000000bffc70000ffedfffb0073ffeaffb1001200010012001fffec0063ffc5fff8ffc100140000000a00b300630027009efffbffa500000000000b0013ffb0ffc500000000000700390000006100120075000d0000, 1024'h001f001b00000000ffe600000010fffbffbeffa4001a003000240046ffd8fff00039ffe1001a0004ffd80000000affaf0000ffe6ff95003cfff0ffe60015004400360008fff100540029ffe20005001d0000ffe4000d008d001400180005ffd4000000000024ffe0ffb4ffb000000000000bfffd000000600030ffc3ffed0000, 1024'hfff1000c00000000fff300000005ffe9ffe9ffb8fffa00090049ffe0ffe30003004200770035fff5ffcb0000000cffdb0000fff7ff8effe10004001f0014004c001cffcc0013000a004affe50047fff30000ffd6ff90003ffffdff9200110006000000000013ffb4000afffb000000000003ffcd000000100025ff74ffdc0000, 1024'hffdcfffc0000000000090000fff2000a001efff6ffccffcb0037ffae0001001600230083002affbeffe700000001fffb0000000dfff3ffc10003003b00130031ffeeffa60024ffef000cfff70046ffd30000ffebff92ffd8fff4ff7b0018000700000000fff4ffc80035003100000000fff5ffdf0000ffce0001ffb0ffec0000, 1024'hfff4fffc0000000000140000ffef003300210037ffbaffd100270003fff900150014000a0023ffbe001700000013fffa000000070065fffdffeb0025000afff5ffebffe10003000fffda0002000afff200000005ffd5ffcffffeffd90009ffe000000000ffebfffa0002000400000000fff7001a0000ffd6fff50005ffff0000, 1024'h001500080000000000020000fff9002bffef0030fff10001001e002effe00007000dffc9000bfff3000900000012ffe30000fff500340024ffe4ffe9fffeffdf00090023ffe600250003ffecffdf00150000fffd000f0017000c0017fff9ffd700000000fff50011ffc7ffd0000000000004002200000012000d000000070000, 1024'h000a000600000000fff2000000030003ffdf000200470026fff1ffd1ffea0007000d000bffd90018ffea00000002ffd70000fff3ffd0001c0003ffd8fff9fff8002b0009ffe3001a0051fff5fff900160000fffd002c003100030003fff9fffb00000000fff20007ffee000500000000000a00060000000c000effe600040000, 1024'hfff3fffa00000000fffe00000001ffd4fffcfff20042000bffc5ffb600050005ffe8002cffce000dffdc0000ffea000900000009ffd7000b0017fffcfffc0014fff8ffcdfff5fffa0019002b001300060000001100260020fff1fffd000a001b00000000fffaffdf001f005300000000fffefff10000ffceffec000200000000, 1024'hffeffff100000000001300000005ffed000affe20007fffbffddffea0007000c00010008fff6fff1fff80000fff2fffc0000000fffe400090017000100050018fffaffe30015fffcfff70000000fffe40000001e002affffffeb000f0018fffd00000000000bfff80012001600000000fffcffe800000006ffdd0014ffff0000, 1024'hffe8fff800000000001900000012000700180006ffe90008ffe2fffcfff800240018ffeefff8ffe3001700000004ffdf000000080020001e000cfff60009fff400200001001400100029fff10016ffdb0000001a0038fff3ffee001f0015ffeb00000000001300020005fff1000000000003ffe90000fff5ffe0002000040000, 1024'hffe7fff800000000000e00000006fffefffc0028002c0008ffbcffe4ffcc00210010ffeaffdbfffefffd00000030000100000001000900250016ffe9000affd200030003ffe50000001d0006fff8001200000015004a002effec0036000dffde00000000002bfff0000f0032000000000007ffff0000ffd7ffd9001bffed0000, 1024'hffe7fffd0000000000180000fff9ffd2ffffffb8000efff6ffcf000b00180015ffdafff3fffd0003ffe20000ffd7000200000014ffc2000700180013000f003effddffdb0011ffefffc60011000bfff200000019002c0018ffeb001c0021000800000000004cfff0fffd0020000000000004ffeb00000009ffcd0012ffed0000, 1024'hffdf00020000000000260000000cfffa000effe3ffc8001d0036004a001300210018fff1003e000600180000fff2ffe30000000200070013000500220009001100170020001efffefff3ffce0001ffe40000fffdffddffe9ffebfffd001efff50000000000540027ffe2ffaf00000000000effe900000036ffdaffdffff80000, 1024'hffd4000f00000000001400000013fffc00050024ffda0011003c0022ffeb00270016000d002e000100040000000ffffb0000fff90028000efffc00180009ffe9000300170006fffe0012ffe20003fffd0000ffd1ffc50006fff2ffe40017fffd00000000005efffdfff2ffda000000000013ffee0000ffedfff3ffc7ffe90000, 1024'hffd300130000000000060000000700040002fffeffeffff70018fffaffed0026001400160017ffecfff500000008ffed0000fffbfffcffffffff00150019000ffff8fff1000800060001ffed0011fff70000ffccffe6000c0000ffe20019fff5000000000064ffeb00010000000000000012fff40000fff0fff5ffdfffdf0000, 1024'hffd3001300000000000700000003000a0005fffdffe8fff300190003ffed00260017000e001cffe7fffc0000000affea0000fffb00050001fffd0019001b0011fff6fff10006000afff7ffee0010fff80000ffceffe700060002ffe70019ffef000000000066ffedfffffffc000000000012fffb0000fff4fff2ffe8ffde0000, 1024'hffe0000d0000000000060000ffd10018fffd000affe1ffdd00270017ffeb001f0009fff50024ffef00070000000dffdd0000fff90013ffd1fff0001400130003ffd6fffeffd500150006fff0000300230000ffe1ffe9fffd0003fff40008fff400000000004effeeffefffee00000000000000250000ffedffef0000ffdb0000, 1024'hffee000500000000000a0000000bffee0003ffe2fff3000f000d0000002c000dfff00011000dfffbfff50000ffe7000a00000003fff5000300040020000b0017ffffffec0012fffdffe7fffe0004fff50000fff2ffdffff9fff6ffe1000e001300000000002c000c0006fffd000000000000fff30000fffafffaffe400060000, 1024'hfff200090000000000100000ffee0003fffe0015fff00010002b002800060012fffdfff900220019001100000000fff70000fffc0021fff4fff600130009ffeffffa0024ffeafffb0001fff7fff200170000ffedffd3ffe7fffcfff1fffc000900000000002b001dffe5ffe2000000000009001700000000fffeffe700050000, 1024'hfff5000f00000000000400000015ffe5000000130005001e000b0010000c0004ffebffff00020029ffff0000ffee001c0000fffb000b000b000000060002ffed00020021000affe2fffb0004fff6fffc0000ffddffe3fff30002fff7fffa001f00000000002d0014fff7fffa000000000010fff10000fff90008ffe5000b0000, 1024'hffe9001500000000fffc00000022ffeafffffff80008001a0008fffb00190001ffef0006fffd0013fff90000ffeb001b0000fff8fff400110008000f000e00020005000a001dffecffe0fff7fff5ffed0000ffcaffeafff40006fff100040016000000000047001a0008fffb000000000011ffeb0000000a0009ffeb00060000, 1024'hffdd001c00000000fffd0000001bfffffffffffcfffa000b001efffe0004000f0005000d000e0002fffb0000fffc00040000fff4fffd000d000100170019000a000600030015fffcffebffed0000fff30000ffbaffdefffc0008ffe5000b000400000000005d000b0002fff1000000000015fff500000005000bffe1fff60000, 1024'hffd8002000000000fffb00000015000400020004ffee0004001e0008fff3001a000e000a0015ffffffff00000008fffb0000fff200090007fffa0017001a000600060006000cfffffffffff1000dfff90000ffb6ffd90004000dffe6000affff00000000006afff7fffefff1000000000019fff70000fff2000bffdfffe60000, 1024'hffde001f00000000fff60000fff40011ffec00090000ffeb002cfff2fff50018fff8000d0013fff6ffe60000fffefff90000fff2ffefffeafff3001100170009ffdefff8fff70001ffe0ffe4fff1000d0000ffb1ffd700080011ffd2000afffa0000000000680002fff1ffff00000000001300110000ffff0008ffd5ffde0000, 1024'hffe0001800000000fffd0000ffc70022ffcbfffd0030ffec005dffc100090016ffe60043001cfff7ffc10000ffebffdd0000fff4ffbeffddfff600270012002bffc9ffd3ffd6000cffbbffcdffce002e0000ffbcffb6000c0008ff960017fff00000000000510029ffdc000f00000000000c003b0000001ffffaff9fffe30000, 1024'hffd500050000000000150000ffb50006ffc8fff8004a0016008bffb0001a001fffed00930035001dffb40000ffe4ffd20000fffbffadffdd0005004efffd003effe0ffc1ffbb0004ffeaffd2ffd9004a0000ffe2ff710016ffe3ff5c0025000700000000002f002bffdc001900000000000500340000000cffe0ff50ffeb0000, 1024'hffc5ffea0000000000320000ffcdffc80004ffff0018002f006effda0025002bfff900ab00440042ffe20000ffebfff200000011ffe4ffc7001a0063ffe7002b0002ffd9ffccffd800460001001a00380000001cff58fff9ffbaff700025003d000000000011fffc0009002000000000fff9ffec0000ffbbffc2ff5dfff40000, 1024'hffccffd300000000003c0000fff4ffbb004f002affc000040004001700170026fff6004700290033003100000005003800000025004cffb10021003affe1ffdefff60012ffffffa800540026003bfffb00000047ffafffb3ffb9ffe60011004d00000000fff9ffd90042001f00000000ffecffb80000ff86ffb3fff200000000, 1024'hffedffd000000000002600000009fff400620045ffafffc6ff8d0027fff70010fff0ffb5ffe4ffff006100000024005100000025007effc5001bffeafff3ffa0ffdf003a001dffae000c00240017ffd20000004f0057ff92ffe10075fffb001400000000ffe7ffeb0053001f00000000ffe9ffd00000ffabffbc00a800120000, 1024'h0019ffe700000000000600000010002e00310027ffd3ffb0ff6c002ffff0fff6ffdfff4dffbbffcc004700000012003200000015006200110003ffb60005ffb6ffd0002f0023fff1ffa10010ffd9ffcd0000003600c8ffc1001100b8fff7ffd000000000ffe9000e0019000500000000fff2000e0000000bffde00ec001e0000, 1024'h002f000500000000ffef0000000b0049ffdeffef0013ffecffc20036ffe4ffee0004ff60ffd4ffd5000d0000000cffdc0000fff400020056ffedffb4000dfff20000002300020043ffa7ffddffb7fffa0000000a00a8002c00270089ffffffa200000000fffe002cffc2ffc6000000000005003c0000006f000a007c00140000, 1024'h001a001500000000ffea0000000c0010ffbfffbf002e003100200022ffe6fff9002bffe90009fffeffd800000005ffb30000ffe8ffae004dfff0ffe8000a00350032fffdffeb00540012ffe0ffef001e0000ffea001900770014000d000bffcd000000000016fffdffb7ffc400000000000e0015000000550023ffcbfff60000, 1024'hfff4001200000000fff700000017ffddffe7ffbcfff9002800460009fff50009003500550033fffeffd00000fffbffd60000fff6ffb0000efffb001e000c004c002effda001000210042fff50038fffb0000ffd9ffa10053fffcffab00150008000000000021ffc1ffecffe700000000000affcb000000090022ff7cffe60000, 1024'hffd8000a00000000000400000020fff80015ffebffc6fff7003dffe3fff00018003e00660037ffd3ffed0000000efffb00000000ffedfff10002002e001700290017ffcf0039fff90026ffeb0048ffc80000ffcfff920000fff9ff9600190002000000000025ffc300220003000000000009ffbe0000ffe80013ff9affe50000, 1024'hffcf0006000000000007000000100020001f0018ffd3ffd60014ffbfffd60023004200470016ffb7ffff00000029fff80000ffff0017fff70004001f00240003ffffffc800240001000effeb0035ffcf0000ffd3ffd1ffeafffeffbc0019ffe000000000002affd000340024000000000006ffe80000ffd7fffdffdeffe60000, 1024'hffdb00020000000000090000ffeb0022000a000dffeeffc6fffbffd7ffcd001f0026001c000cffbcfff400000029ffed00000003000cfff7000200180026000effd7ffc3fff60011ffe6fffe001afffd0000ffedffff000dfffeffeb001bffd0000000000032ffc9001a003300000000fffd00110000ffdaffe90006ffdf0000, 1024'hfff2ffff0000000000120000ffd30019fffcffdeffd4ffcf00250028ffe700140016fffe0037ffd3fff60000000bffd800000007fff5ffebfff50021001a0033ffd4ffdcfff00019ffd3fff2000e000b00000006ffe60013fffdfff2001affd600000000002affdaffe6fff300000000fff9001900000012ffe8fff5ffe20000, 1024'hfffbfffc0000000000130000ffde0017fffafff5ffccfff80055003bffee001000270012004dfffb000700000013ffd80000ffffffffffe4fff0001e000200150001000dfff1000b000effd9000a000f00000006ffb20002fff8ffd6000bffe800000000000bfffcffd9ffc400000000ffff000b00000020fffaffc0ffeb0000, 1024'hfffbfffc0000000000090000fff700040008001cffe80003002ffff500000010000b002c0019ffff00010000fffbfff3000000020014ffe8fff70009fff2fff5000b0004fffffff80032fff30010fffa00000000ffc8ffe8fff7ffc80000000f00000000ffe8fffefffbfff4000000000000fff30000ffec0002ffcbffff0000, 1024'hfff8fff800000000000200000007fffc0009002d001f000bffe2ffcbffff0008fff90018ffdf000400010000000b001400000003001c000a000bfffbfff6ffdb0006fff8fff7fff200120012fffb00040000000b000dfff4fff6fffafffd000800000000ffe90008001c003200000000000000000000ffd0fff5000600080000, 1024'hfff6fff60000000000070000000fffe4fffffff90033000dffc1ffd300090005ffe90004ffd60011fff00000fff6001b0000000affe20017001bfff4fffbfffdfffcfff1000affe8fff50012fffcfff50000001600360007fff200180009000c000000000009000600190035000000000005fff20000fff3ffe8001500020000, 1024'hffeefffc00000000001300000010ffe5000fffe0fffb0012ffe000140027000effe6ffe9fffa001000070000ffe1000a0000000afffe0015000e000dfffd0012000600010019fff1ffe600070003ffe9000000150020fff2fff3001d0010000f00000000002700140000fffb000000000006ffed00000002ffdf001a00020000, 1024'hffeffffc00000000000e0000fff2000bffe90022002600170007ffe3fffe001efff3fff8fff10010fff900000003ffec0000fffcffeffffa000affe8fffbffd200010022ffe5fffc001affcfffd100140000fffe001cfffffff000020009fff80000000000290039fff0fff3000000000006000b00000011ffe4ffee00000000, 1024'hffdcfff60000000000150000ffdfffebffe10000006e0008fff4ff9b0010001affcc004affdf001fffc00000ffe8000b0000000cffbc00080021001cfffc001bffd4ffc5ffd6ffe5ffd00008ffda002b0000000a0005001cffdfffd20023000a00000000002a0015000a0061000000000005001a0000ffe7ffc7ffd0fff90000, 1024'hffd0fff60000000000350000000dffc40018ffbfffe900320021002e00460029ffe80027002e0024fffc0000ffbefff500000017fff4001c00170044fff600460015ffef001effedfff200000016ffe80000001fffd3fff5ffd1ffe3003400250000000000480010ffeeffe4000000000009ffcf0000ffffffbdffcc00060000, 1024'hffcd000000000000002b00000025fff50011002cffb80029004c0058fffe00360017fff40047001300190000000e000b0000ffff00440019fffd001afff6ffd200170041001affef001affcbfff6ffed0000ffe8ffbbfff9ffdffff1002100000000000000660015ffe2ffaa000000000015ffd10000fff8ffe0ffbdfff10000, 1024'hffc8000f00000000000e0000000900050004000effeefffc001c0002ffec003100120010001cfff5fffb0000000ffff60000fffc000a0002000200170012fffefff6ffff0004fffd0000ffe50006fffc0000ffcdffe50008fff8ffe7001ffff4000000000077fff50000fffb000000000016fff30000ffeaffe7ffddffda0000, 1024'hffc8001100000000000c0000000200040007fff8ffedfff500130002fff1003000110010001bffeefffb00000006ffea0000fffefffffffe0002001c00190014fff2fff200050003fff6ffed000ffff90000ffcfffed0006fffdffea0021fff300000000007bffed00010001000000000015fff60000ffefffe4ffeaffd80000, 1024'hffd8000b00000000000c0000ffc8001600020009ffd4ffd7002a0028fff200260002ffea002dffef000e0000000affde0000fffc001effc6ffef001b00120003ffc90001ffcf0015fffdfff0000000290000ffe4ffe8fff6fffffffb000dfff7000000000061ffefffedffe700000000fffe00290000ffe7ffe2000bffd50000, 1024'hffe1000000000000000900000014fff50008ffe0fff5fff6fff2ffe500090010000a001d0002ffdeffec00000009001200000005ffeb00060010001f001d0019fff5ffce00170001ffe800010018ffed0000fff0fff40016fff1ffec001bfffb000000000034ffdd0024001d00000000fff8ffe80000ffe3fff7fff4fffc0000, 1024'hfff300020000000000170000ffcc0020fffefff1ffd5ffd9002d0021fffd001e0005fffb0031ffe400030000ffffffd7000000070006ffd5fff1001a001b0019ffdbfff9ffea000dffe7ffe90002000e0000fffeffdfffedfffcffe6000effea000000000028fffeffe0ffe600000000fffa00230000000dfff2fff4fff90000, 1024'hfffd00050000000000130000fff9000900020023fff2001a00270027000000130005fffa001b001e001200000003fff70000fffd002a000afff4000dfffeffe80011002afff0fff7000efff6fff3000f0000fffcffd8ffedfffcfff1fffb000100000000000f0021ffddffe100000000000b000e0000fffffffeffdd000c0000, 1024'hfff5000c0000000000020000002bffd40002001300140038fff5000b00180004ffe6fffdfff0003700000000ffed00290000fffb000a001e0008fffffff8ffe3001a00280011ffdf000f000cfff5fff90000ffe6fff2fffffffc0003fff9002a00000000002900190000ffff000000000012ffdd0000ffec0007ffe600100000, 1024'hffe3001200000000fffc0000002affdf0002fff60016001cffecfff4001d0005ffe2fffeffee0024fffa0000ffea002c0000fffbffed0011001000070007fffc000500110022ffdbffe60000fff7ffea0000ffd00001fff20003000200030022000000000052001a00130009000000000017ffe30000ffff0002fffaffff0000, 1024'hffd9001800000000fffe00000007fffffff1fffb001400030015ffe700170012ffdf00090002000fffea0000ffe700110000fff7ffe6000000040013000d0008ffe7ffff000fffe9ffc6ffe4ffe5fff80000ffbfffecffee000affe1000e000b0000000000680027fffc0002000000000019000900000010fffaffe4ffef0000, 1024'hffd200100000000000040000ffcd000cffcd000300470009004bffba000b001bffe7004800140015ffca0000fff3ffea0000fff3ffbaffe50007002700090014ffd3ffe3ffcffffbffd2ffcfffcb00350000ffc8ffbd0008fffaffa50017fffd0000000000600036ffed0019000000000011003500000018ffe6ff9fffe00000, 1024'hffc2fff500000000001f0000ffb4ffd8ffecffed00480017004affb200170024ffee00940025003affd50000ffeeffe300000008ffb3ffba001f004efffb0032ffdcffcbffb6ffe3001efffc0004004a00000004ff92fffdffcfff8c0020002d00000000003a000a0011003e00000000ffff00190000ffdbffbfff8affe00000, 1024'hffc3ffd200000000003a0000ffd6ffb50040000cffe8ffff0002fff000150027fff0006900220039001d0000fffb001d000000260016ff9d002c0041ffe9fffdffe2fff6ffe7ffab00500026003c000f00000047ffb4ffbbffb7ffd8001a004f000000000007ffd60049003c00000000ffebffcc0000ff93ffa2ffebfff60000, 1024'hffe3ffc900000000003400000005ffe6006a0038ff9dffc3ff9f002c000c0019ffe2ffccfff8fffb005a0000000f0053000000300081ffbe001d0000ffecffb6ffd300280027ffa6000000290022ffc90000005b003cff86ffd4005d000a002300000000ffeaffe50053002000000000ffe7ffc50000ffa0ffac009500100000, 1024'h0014ffe200000000001200000014003a003a003affb7ffbbff83004dfff10002ffedff42ffd1ffcd005b0000001b002d000000140086001afffcffbcfffdffa4ffdf00460025fff3ffac0001ffd5ffc90000003d00b8ffb2000c00b7fffaffc800000000ffeb001d000cffe500000000fff5000c0000000dffd600e3001f0000, 1024'h0030000800000000ffee0000000c004dffe0000a000fffefffbc003bffddfff60001ff4bffc9ffd100160000000cffd20000fff2001f0058ffe6ffa3000bffdb00050033fff50050ffc3ffdfffb100010000000700be002d00280099fffaffa300000000ffff002dffb9ffbe000000000004003b0000005d000b008c001a0000, 1024'h0021001900000000ffe300000008001affb6ffcb004400280005001affd7fff70022ffccffeffff5ffd400000008ffad0000ffe5ffb5005cffedffd30011002b0028fffcffdb0065000affeaffdf002a0000ffe800470089001b002c0007ffbf000000000015fff8ffb0ffd200000000000d0026000000520025ffedfffc0000, 1024'hfff9001100000000fff300000014ffdfffdcffa50012002800330001ffe300060041004f00260000ffc800000001ffc30000fff4ff8e001a000100110012005b0034ffd30007002e004ffff4003c00020000ffe0ffc30070fffdffc10018fffa000000000021ffb4ffeaffec00000000000affd10000001c0020ff87ffe40000, 1024'hffd500030000000000070000001fffec0019ffd4ffc3fff20032ffe1ffed001b00440074003affd4ffe70000000efff900000006ffd8ffe9000800310015003b0016ffc1003efff40034fff2005fffc20000ffddff94000bfff3ff9600210007000000000022ffa9002b000c000000000006ffb10000ffe0000cff98ffdc0000, 1024'hffcc000200000000000d00000023001b002d000effb2ffd50016ffddffe0002600450044002bffb100060000002c000c000000060023ffff0004002e001e000c0005ffcb0042fff0fff3ffec003fffb80000ffdaffbdffe2fffdffb90021ffde000000000032ffcb0036001b00000000000bffcf0000ffd6fff9ffd7ffdc0000, 1024'hffcf000d00000000000900000021001f0017000bffd0ffe70003fff0ffdb002b003a00110019ffbe000500000029fffa0000fffd001b001c00020018002400020008ffe2002c0006ffebffe60021ffce0000ffd2fff0fffd0004ffe6001fffd0000000000058ffe20019000a000000000014ffe70000ffeefff6fff0ffdc0000, 1024'hffcf00160000000000070000000f00150008fffbffe5fff00005fff8ffd8002f003400040012ffcefffe00000019ffd90000fff8000200130000000e002a000f0006ffe9000e001b0009ffe6001dffe90000ffcb000600150003fff5001dffd8000000000070ffe00004fffe000000000012fff20000fff7fff3fff4ffdc0000, 1024'hffce00100000000000080000fff000100003fffffff5ffe20001ffefffc5002d0030000e000effd6fffb00000024ffcf0000fffafff7fff30004000b002f000cffecffe4ffeb001d001cfff0001e00080000ffd500090020fffdfffd001bffdc00000000006bffcb000c001100000000000700040000ffe7ffe9ffffffd80000, 1024'hffd7000100000000000e0000ffd5000c0007ffeaffeaffbefffffff8ffc9002200200016001cffd4fff40000001fffe000000008ffe8ffd200060017002a0024ffc6ffd0ffe9000afff7fffe0025000c0000fff1fffd0017fff7fffa001fffe000000000004fffb60012002300000000fffb000c0000ffe8ffde000affd40000, 1024'hffe9fff50000000000180000ffcf001d0010ffe2ffc2ffc0001d0018ffe7001d001e000b0037ffcf00070000000dffd80000000efffbffcbfffb001c00170027ffd3ffe2fffd0006ffedffe90020fff60000000effe9ffedfff8ffee001bffdf000000000020ffd7fffdfff500000000fff6000d0000000affdf0005ffe30000, 1024'hfffbfff50000000000150000ffe4002000100015ffc4ffe70027002cffee0015001efff90031ffe2001a00000018ffe6000000060034ffeefff000110002fff7fff40007fff6000cfffefff00008000200000014ffdfffe8fffafff60009ffe300000000fffbfffbffefffe200000000fffb00130000fffeffeefffdfff40000, 1024'h0009fffa00000000000600000001000c0005001efff0000700020011fff4000a000effef0002fffb00100000000efff30000000000210003fff7fff0fffaffe2000f0019fff600090022fffbfffd00040000000d0009fffefffd000bfffbfff800000000ffed0004fff4ffef00000000fffdfffd0000fff60000000400070000, 1024'h0001fff800000000fffd0000000ffffbfff9000f0035000fffcdffcdfff80006fff50005ffd20011fff500000007001000000002ffec00140010ffe4fff8ffe6000b0004fffeffee00160007fff7fffe0000000b0030000bfffc0011ffff000400000000fff5000400130029000000000006fff90000fff1fffb000b00080000, 1024'hfff6fff800000000000700000009ffe8fffeffe000270003ffd6ffe000230004ffd70009ffe3000fffe40000ffde001e0000000cffda00140011000afff8001dffeeffe00010ffe8ffcc0011fff6fff50000000e001f0008fff700040013000f0000000000120006000c002e000000000003fff70000fffbffe5000900050000, 1024'hffecffef0000000000140000ffef0002fff3fff00020001a0013ffe5001000160007001e00040013fff90000fffeffe700000003ffd0fff300130006fffa000200090005ffedfffd0014ffd5ffea000f0000001000010000ffe7ffed0017fffd0000000000180026fffffff500000000fffc00000000001cffdbffe100030000, 1024'hffd2ffdf00000000001e0000ffeeffee0002000c00480000ffefff90ffef00270001006dffe90011ffdc0000000d000600000015ffc9ffeb002c0010fff80004fff0ffd0ffe9ffd8002bfffb000a000c0000001efffc000cffd0ffcd002a000a000000000008ffe60034005b00000000fffbffe90000ffccffc3ffd0fffb0000, 1024'hffc5ffe000000000003500000023ffd0003affcdffd8fff5ffd100030030002fffea002c0011fff4fffb0000ffe100320000002b000f001d00230040fffa003cfff5ffc10047ffccffc300210032ffbc00000035fffcffecffd1fff700430010000000000031ffd4002c0036000000000004ffb70000ffc2ffb00007fffb0000, 1024'hffcdfff00000000000310000002e000e001d0000ffa3001c002000670002003c0035ffcf004afff4002d000000210007000000060030002a00060017fffdffe30025003c003afff0fff3ffb7fffcffc900000008ffeeffedffe40016002dffd600000000006d001fffecffa2000000000016ffc900000024ffccffe9ffe70000, 1024'hffc2000a0000000000170000000900080004000effe600020020000fffea003d001a00070026fff3000000000011ffed0000fffd000c0007000200140010fff8fff8000a0006ffff0005ffd80002fff70000ffd3ffea0006fff3ffec0026ffed000000000085fffbfff8ffed000000000019ffef0000fff5ffdbffdaffd60000, 1024'hffbd001000000000001200000002ffff0007fff8fff0fff90011fffdfff1003b00100015001cffecfff800000003ffe500000000000000040005001e001b0014ffeeffed00050005fff7ffec0010fff70000ffcefff00007fff8ffe9002afff300000000008dffed00020006000000000019fff60000ffeaffd9ffe7ffd50000, 1024'hffd1000a0000000000130000ffbf001400040006ffc9ffd5002d003afff4002e0002ffdf0038ffed001300000008ffd70000fffd0029ffc4ffec002200140006ffbf0001ffc6001cfffafff4000200300000ffe8ffe9fff5fffb00020011fff7000000000072ffebffe6ffe100000000fffd00300000ffe2ffd70012ffcf0000, 1024'hffcf00090000000000070000002bfffd000bffeb00000004ffebffd0fff40019002a0020fff6ffd9ffef0000001b00080000fffaffeb00230017001e002700150015ffcb001b000e0008fff60022ffe40000ffde00070027fff1ffef001effeb00000000004effd8002c001d00000000ffffffd80000ffdefff7ffeefff40000, 1024'hffe000030000000000130000ffb90024fffdffefffe0ffac00230008ffca002300110010002bffceffee0000001bffcf00000008ffecffbefffa0021002e002dffb8ffd3ffd10012ffe9ffef001100240000fff3ffea001cfff7ffec001fffd4000000000047ffbcfff6000e00000000fff000200000fff0ffdffffdffdd0000, 1024'hfff7fffb00000000001b0000ffd5002a000afff0ffc2ffd4003e002efff400210014000a003effdf000800000006ffce0000000c000effdcffee002000100025fff1fff9fff7000bfff3ffe1000c00040000000bffd0fff4fff8ffde0018ffdd000000000011fff3ffddffd800000000fffb001000000010ffecffe5fff80000, 1024'hfffc00010000000000110000001c000c000e0027ffd80026002400320005001b0016fff7001d000c001a0000000effff0000fffd00410021fff00009fff6ffdd0030002e000bffff0021fff1fffdfff80000fffcffd6fff7fffafff10002fffb0000000000090017ffe5ffd100000000000dffee0000fff10005ffd7000d0000, 1024'hfff5000c00000000fffc00000026fff0fff2001e00220026fff5fff3000b000fffe8fff8ffe90027fff00000fff600270000fff8000000220001fff0fff4ffdc000d0020000bffe60006fffdffe8fffc0000ffdb0003000b0003fffafffe001800000000002f0017fff80007000000000017ffee0000fff0000cffe100030000, 1024'hffde000700000000fffc0000fff5ffebffe0ffeb005a001afff6ffb6001e000dffd6002effe40035ffd50000ffe900170000fffbffadfff80018000ffffc000effeafff0ffefffdbffdffff3ffdf00180000ffe0fffb0007fffdffdb000d001a00000000004a0027000c0034000000000012001000000005ffebffd6fff00000, 1024'hffcbffef0000000000160000ffd1ffce0003ffe70045001cfffcffb40029001effe3005efff7003dfff50000ffeafffa0000000cffbeffba00290028fff90011ffecffeaffd2ffd5002800060004002b00000010ffe0ffe1ffd7ffcf0013003a0000000000350017002f004000000000fffd00010000ffdaffbfffdefff20000, 1024'hffd5ffdb00000000002e0000ffdbffd600360021fff9ffdcffd4ffd5001c0023ffcb0022ffed001000160000ffde001f00000026002bffb50020000ffff2ffe7ffbefff2fff2ffc4001200230011fffb000000340017ffacffcd00080017003d000000000005fff2003c004400000000ffebffee0000ffaaffad003e000f0000, 1024'hfff9ffe10000000000280000fff20020002e0034ffd4ffccffb7001b0004001affe0ff9affe1ffd500350000fff400090000001c0072000e0003ffe0fffcffcaffcf001100070002ffc90007ffe4ffdf0000003f0080ffbafff0006a0014ffe400000000fff000150002ffff00000000fff0001a0000ffecffc0009b00240000, 1024'h001ffffd00000000000c000000020039ffed0019fff40000ffd9005fffe1000d0007ff5fffefffd8001d0000000dffcd0000fffb004c0061ffe5ffc30002ffda0004002fffe90052ffd5fff0ffc1000c000000250090002e000c00870008ffac000000000001001effadffb9000000000002003800000037fff0006c00140000, 1024'h0023001400000000fff60000000b000effc2ffd10012002a001b0058ffd800010024ffb20010fff7ffe20000ffffffac0000ffebffd3005bffe4ffd50009002100240017ffe700600011ffe3ffe5001e0000fff60036008100100038000cffc500000000001efff5ff9affa800000000000c0015000000580019ffe7fffb0000, 1024'hfffc001300000000fff600000013ffedffd6ffb10001002a004c0017ffe200070045003f0037fff8ffcd00000005ffbe0000fff0ff9e0020fff800100012004e002fffe200080036003dffe1002b00020000ffd8ffb7006a0001ffc00019ffee000000000029ffc7ffd9ffd000000000000cffdd000000300023ff80ffe40000, 1024'hffd400080000000000040000001cfff1000dffd4ffcffffc0047ffd8ffe5001c005200850040ffd3ffde00000013ffe900000000ffcbffef00060034001a0041001effbc00330002003effe9005cffcd0000ffd0ff84001afff4ff8300230000000000000027ffab00230008000000000008ffb70000ffe90013ff7dffdb0000, 1024'hffc3000500000000000e000000210013002b000affb8ffd6001cffc6ffde002d0048005e002bffaefffa000000230004000000070018fffb00070031002100170007ffba0043fff3000bffee0050ffb20000ffd4ffb3ffe5fff9ffa20025ffe7000000000033ffbc0039002500000000000cffc80000ffc9fffdffc3ffdb0000, 1024'hffc9000c00000000000d0000001b0024001f0017ffccffddfffcffe9ffd20031003f00120017ffb600090000002efff60000fffe002d001d0001001c002500000004ffd800270009fff1ffef002affce0000ffd9fff7fff90002ffe8001fffcb000000000054ffd8001d0017000000000013ffed0000ffdcffeefffaffd60000, 1024'hffd0001600000000000800000016000e0007fffdffe6fff6fff70008ffd40031002cfff40011ffd600000000001effdf0000fff90007002000010009002500080007fff4001200140001ffec001affe90000ffd30011001c00040009001dffd600000000007affe30000fffe00000000001afff10000fff6ffedfffbffd10000, 1024'hffca001900000000000700000016ffff0002ffeffff20002fffd0004ffe30033002000000010ffebfff900000011ffe10000fff8ffee00120005000d002400100008fffa000f000a000affe90018fff00000ffc80006001d0001fffe001effea00000000008fffea0001fffc00000000001cffe80000fff8ffecffebffd10000, 1024'hffc1001a00000000000a0000000cfffe0007fff7ffedfff80008fffeffec0035001200080014ffecfffa00000006ffe90000fffbfff800010005001700250011fff6fff6000b0002fffeffea0014fff20000ffbffff800090000fff10020fff5000000000099ffed0005000100000000001affec0000ffeeffe7ffecffd50000, 1024'hffc0001900000000000b0000fff6000f00050007ffefffe90010fff3ffe10036001800040011ffdeffff00000009ffd80000fff90005fff300010010002d0007ffe9fff3fff800130003ffe2000afffc0000ffbd000200000000fff2001effe900000000008efff00001000000000000001200010000fff1ffe5fffcffdf0000, 1024'hffc7001100000000000c0000ffe0001a0000000cffffffd50007ffe5ffc400310023000a000bffd2fffa0000001cffc90000fffb0003ffef0003000c0032000affd8ffe0ffdd0021000affef000e00120000ffd000130014fffbfffe001effd8000000000072ffd50006001800000000000700180000ffe8ffdf000cffdd0000, 1024'hffd900050000000000120000ffcf00150000ffedffe9ffbf00090000ffc60027001e0007001dffcafff100000014ffc900000006fff3ffe3ffff0012002c0027ffc4ffceffe10020fff5fff8001d000f0000fff1000c001ffff800020024ffd5000000000051ffbbfffc001300000000fffb001b0000fff2ffdb000fffda0000, 1024'hfff0fffd0000000000180000ffd000200007ffe6ffbbffcf002a0039ffde00210029fff50040ffcb000a00000012ffbf00000008000dffe1fff00018001a0026ffe2ffecffed0025fffcffeb001d00070000000dffed0009fff9fffc001affd3000000000026ffd5ffe1ffdb00000000fff700160000000bffe60001ffe20000, 1024'h0004ffff0000000000100000ffe8002400000017ffc5ffeb00380036ffdf00150025fff00034ffe0000c00000017ffd7000000000025fff5ffe800040005fffbfffd000ffff1001b0011ffe30005000700000006ffe00006fffffff20007ffdc000000000001fff4ffd6ffcd00000000fffc000c0000000affffffe6fff20000, 1024'h0002ffff0000000000000000fffb001effee001c0019fffe0017ffd6ffe5000e0013001bfff9fff8ffea0000000dffeb0000fffbffef0009fffcfff1fffafff7000efffafff30009001effe3fff600050000fffaffff0016ffffffde0007ffe900000000ffee0002fff000030000000000030004000000050005ffd5fffd0000, 1024'hffecfff70000000000040000ffffffeffff9fff500390013ffecffc00003000efffc003fffea000bffe100000003000200000006ffdb001200160014fff80017000dffd2fff3fff9000f000f0008000e00000013fffc0023ffeeffe10013000100000000fffefff00016003e000000000002fff70000ffdbffe8ffdbfff70000, 1024'hffe8ffee00000000001800000001ffea000affe60006fffbfffeffd7000a001800070033ffffffeeffe70000ffeafff300000011ffd6fff80014000b00020022fffeffd50012fffe0013fff40012ffe8000000150004000bffdfffe100230005000000000009ffee0013001900000000fff7ffd50000fffbffd9ffe400030000, 1024'hffceffe700000000002300000010000e00180009000bfffbffe6ffafffdb00320037003cfff4ffd3ffff0000001bffe00000000ffffe001f002200010010fffe0016ffd2001600070034ffe60025ffd2000000190028fffdffdbfff30031ffdc00000000000effe4002d0026000000000002ffe20000ffe9ffcdfffd00010000, 1024'hffc6ffee0000000000270000002dffed0024fff2ffebfff7ffb5fffbffe0003d001f000a0000ffd5fff80000001f000e00000017001c004a001b001a000f00130006ffc9002cfff7fff4001c0037ffce000000230030002cffde0020003bffda000000000048ffb30022003e00000000000fffcc0000ffb8ffc00011ffdf0000, 1024'hffcffffa00000000002800000026fff70016ffc7ffba000cffeb004cfff600430033ffd1002fffe100110000000cffe10000000afff00028000c000a00130016001a0010003700030004ffd30023ffc50000000a00240015ffea00290034ffda000000000088ffeffff3ffc9000000000016ffc200000020ffc6ffffffd30000, 1024'hffbb000800000000001f00000007000600070002ffdf000100170013ffe5004600240001002bffec000400000012ffe30000000000030009000800130018fffbfff50009000cffff0003ffd0000affec0000ffd8fff60001fff0fff6002effe6000000000099fffbfffaffe900000000001bffee00000001ffcfffe2ffd10000, 1024'hffb2000f00000000001a00000001fffa0009fff8fff0fffc000dfffbfff1004600130018001fffecfff800000004ffe40000000200000004000a0022001f0011ffebffec00060001fff7ffea0013fff40000ffcffff10004fff1ffe80030fff300000000009fffee0004000b00000000001bfff40000ffe5ffcfffe5ffd10000, 1024'hffcb000a00000000001c0000ffb5000f000a0005ffbcffd0002f004afff80034fffdffd50041ffec001900000002ffd4000000000034ffbdffec002b00170008ffb10001ffc0001cfff2fff8000400340000ffedffe8ffedfff600090014fffb000000000083ffeaffe3ffdd00000000fffa00360000ffddffca001cffcb0000, 1024'hffc0000e00000000000a00000048fff30012ffe2fffc0011ffeeffc3000c002500220029fff4ffe0ffe80000ffff00160000fffbffe10037001a0023001e00200021ffc8003dffff0003ffeb0028ffc30000ffca00040017fff2ffdc002afffd000000000070ffe70030001600000000000effbe0000ffe5fff2ffdafff10000, 1024'hffbe00080000000000120000ffbf002d00000009ffefffb40024ffedffaf0034002e001c0025ffccfff60000002fffc40000fffffffaffcc000100200034001effc0ffd1ffc6001f0004ffe2001300250000ffd8fff7001efff8ffec002affc6000000000072ffb70002001600000000fffb00200000ffe1ffd2ffffffcf0000, 1024'hffd9fffc0000000000170000ffbf00210008ffe2ffc6ffac0027001effcb002b002000170041ffbefff700000020ffc60000000ffffcffc5fff800290027003cffc7ffccffe4001affecfff20022001300000004ffdf001bfff3ffe90029ffc900000000003effb0fff4000600000000fff6000f0000ffedffd8fff9ffd10000, 1024'hfff5fffe00000000001c0000ffef0027000bfff5ffa4ffe300450047fff500240028fffa0050ffcb000c00000011ffd500000007001ffff5ffe90021001000190003000000110014ffeeffd6000fffee00000007ffc5fffafff8ffdd0018ffd100000000001dfffaffd7ffc2000000000001fffb00000018fff3ffd4ffec0000, 1024'hfff4000300000000000f0000fffa0020ffe8002c000600170047fff8ffef001d0017001e0023000bfff100000015fff20000fff500020010fff6000cfff7ffe600100015fff0fffb0011ffceffe7000f0000ffedffc30006fff9ffc20008ffeb0000000000180025ffddffe5000000000010000f00000010ffffffa1fff20000, 1024'hffe0fffa00000000000c0000ffdfffe9ffee000c0051001c0010ffa20016001dffdf005bffea0032ffd70000ffe3fff700000003ffcdffe800130016ffec000afff9ffe2ffd2ffe6002e0000fff8002700000002ffe20003ffe7ffb8000f002800000000001100110009003c00000000000400090000ffd5ffdcffb8fffa0000, 1024'hffe6ffee00000000001f0000ffcfffecfffc00170030fff60007ffb000340021ffb30033ffe3ffffffd90000ffb7fff400000018fffdffe1000d000cffee000bffc9ffcfffddfffbfff00005ffdc00140000001c000effe5ffdaffd10020002400000000fffc001efffc003800000000fff0000e0000ffd5ffc2fff6001a0000, 1024'hfff1ffee00000000002c0000ffe20016fff0001d001e000e0020fffe0009001ffff2fff90006ffedfff30000ffebffd60000000b002a003c0003000dfffb0002ffefffe8ffd90030ffd7fff0ffc9001c0000002a001e0010ffdb00040028ffd900000000fffc002affd0fff900000000fff900300000000dffc7fffd001e0000, 1024'hfff8fffa00000000002800000003fff1ffedffe4ffe9002d003c005effec001f0023fff4003a0001fff00000fffcffc200000002000a004bfff7001500000025001c0000ffed003c001efff20005001500000020ffed005bffdd000c002affde00000000001cffe2ffb5ffba000000000000fff900000015ffe3ffc300030000, 1024'hfff1ffff00000000001b00000010ffecfff8ffd0ffb600170057005dffdd001e0048001d005fffecffef00000011ffd000000001ffe60015fff6001d000b002e001dffff001400210035ffdb0030fff20000fffdffa9004bffe7ffd90027ffe8000000000031ffbfffd4ffb0000000000003ffca0000001bfffeff94ffe50000, 1024'hffd5000000000000001300000019ffff0013ffdeffb1fff6004b000affd800210060005d0057ffcdfff400000027ffed00000003ffe6fff700040033001d002d0017ffd80037ffff0023ffd8004dffc90000ffdfff8a0011fff0ffa20027ffe6000000000033ffb80015ffeb000000000008ffbe000000010005ff90ffdb0000, 1024'hffc1000400000000001300000023000d0028fff8ffb1ffdd0027ffd5ffdb002d00570061003affb0fff900000026fffe000000060005fffb000a00350028001f000affbe004afff4000bffe20054ffad0000ffd2ffa7ffecfff5ffa0002affe3000000000040ffbb0036001600000000000cffc10000ffdffffcffb5ffda0000, 1024'hffbe000c0000000000130000001d00210023000fffc0ffd9000bffdcffd200380049002d0024ffab00030000002cfff2000000010023001400050027002d000b0002ffca00340005fff6ffe6003affbf0000ffd1ffe0fff1fffdffce0028ffce00000000005effd000260018000000000013ffe20000ffdbffeeffe4ffd40000, 1024'hffc5001400000000000f000000130019000e0008ffddffedfffffffeffd0003c003300020019ffcd000100000026ffe10000fffa0015001f00000016002800060002ffea0013000ffffcffea0020ffe50000ffd1000200120001fff80023ffd0000000000080ffde0006000700000000001bfff50000ffe8ffe6fff2ffcc0000, 1024'hffc8001800000000000c0000000c00050003fff5ffeafff90007000cffe0003a001dfffc0018ffe7fff90000000cffdb0000fffafff800100000001000210011fffcfff90008000c0004ffe70015fff40000ffc90003001a0000fffc0023ffe7000000000095ffe7fff8fff800000000001cfff00000fff7ffe3ffebffce0000, 1024'hffc0001800000000000c0000000b00010001fff6fff3000100100001ffed003c0014000b0018fff0fff800000006ffe00000fffafff60007000300140020000dfff9fffc000800060001ffe3000dfff60000ffbffff5000efffeffee0025fff200000000009cfff3fffdfffa00000000001efff20000fff5ffe4ffe3ffd40000, 1024'hffba001800000000000e0000000c00020004fffdfff5ffff0010fff5fff10040001200120015ffeefff700000004ffe50000fffbfffc0006000400180021000bfff5fff600080004ffffffe5000dfff50000ffbafff30007fffcffe60027fff60000000000a1fff50003000300000000001efff30000ffebffe2ffe2ffd60000, 1024'hffb7001800000000001000000003000300010001fff9fffd000ffff9fff10042000a000c0016fff4fff700000004ffe80000fffb000100040003001a00210008ffeafff8ffff0002fff5ffe80007fffd0000ffbbfff40005fffdffea0027fff60000000000a8fff7fffe000600000000001fffff0000ffe7ffdeffe7ffd40000, 1024'hffba00180000000000110000fffb00000001fffcfff5fffe00150003fff1003f000e0009001afff1fffa00000001ffdc0000fffbfffefffc0002001b0026000dffeafffafff7000bfff9ffe6000400040000ffbdfff30008fffbffed0026fff40000000000a7fff8fff9ffff000000000019fffd0000ffefffdbffe9ffda0000, 1024'hffba00160000000000130000fff9000600040000fff0ffef0019fff7ffdd003c00200010001affdffffa00000007ffd30000fffcfffefff9000500140030000effe5ffeffff800160007ffe2000ffffc0000ffbbfffa0009fff7ffed0029ffec00000000009affe50001ffff000000000012fffb0000fff3ffdffff0ffe10000, 1024'hffba000d0000000000140000ffe300160005fffcffecffcf0011ffedffbf00380032001a001fffccfff600000023ffcf0000fffffffaffeb0007001b00380018ffd2ffd4ffea001b0005ffe8002000050000ffcefffd0019fff6fff1002cffd4000000000083ffbf000c0015000000000006000c0000ffe5ffdbfffcffd60000, 1024'hffd100040000000000190000ffc100230001ffe6ffc9ffad00290010ffca003000250010003effb7ffef00000018ffc400000009fff5ffcefff7002600310037ffb7ffc5ffe60021ffe0ffe80020000b0000ffeeffe80016fff8ffe5002cffca00000000005effb9fff2000500000000fff9001c0000fff7ffd9fff8ffcd0000, 1024'hffe9fffc00000000001d0000ffba0034fff7fff8ffc4ffcd0058002cffd90027002b00110058ffd3fffe0000001cffbd000000040003ffd5ffec002800140025ffdaffecffde001cfff0ffd1000a001700000007ffbf0002fff8ffcf001cffc8000000000029ffedffd2ffd700000000fffd002a00000019ffe3ffcdffd50000, 1024'hffeffff50000000000170000ffd70011fffb001bfff2000000470001ffe7001d001d003600340008fffc00000012ffdb000000020004ffe5fff9001afff2000400040000ffdffffe0033ffe4000a001800000013ffbafffdffeeffc1000bfff400000000fffaffffffe7fff200000000000300090000fff8ffe8ffafffe60000, 1024'hffedfff00000000000110000fff7ffe80008001b0014000a0003ffcf000f0014ffe9003afff8000affee0000ffee00090000000c0005fff5000c000dffebfff8fffcffeafffaffe8001900090002000000000019ffe9fff4ffe5ffd5000e001800000000ffec0001000f002b00000000fffeffea0000ffd2ffdeffda00010000, 1024'hffe3ffee0000000000180000001bffe9000b000600200014ffe6ffce0001001100080029fff1fffafff30000000200130000000efff4002a0024000efffb0001000dffe20016ffecfff5fffe0000ffe80000001900120004ffddfff9001ffff900000000000c00070021002e000000000004ffdb0000fff5ffd3fff000030000, 1024'hffcafff800000000002300000037ffe5001affdffff80015ffe0ffddfffe002e00210022fffbffe5fff50000fff5fff60000000effeb003a0024000c0010001a0025ffdb0042fffb0018ffeb002dffb4000000080024000cffddffff0035fff400000000003fffe8001d000a00000000000dffb90000fff9ffd4fff2fffd0000, 1024'hffb900000000000000230000002cffff00190000ffe70008ffdffffaffdc004900330007000cffd8000300000029fff0000000060014003a00180015001afffc001affe9002300040013ffec0027ffd70000fffa001e0021ffe200100036ffd500000000007affdd0018000e000000000017ffd50000ffd6ffc9fff8ffd40000, 1024'hffbc00090000000000220000000ffff50010ffe8ffddfff8ffeb0019ffe4004d001ffff2001bffdffffc0000000cffdf00000008fff80016000d001300210014fff8fff2001400050002ffea0020ffe50000ffeb001b001effeb00110035ffe30000000000a4ffddffff0000000000000018ffdc0000ffedffc3fffaffc90000, 1024'hffb2000b0000000000220000000200020007fff2ffecfffd00090007ffe7004e001f00040021ffecfffe0000000bffd800000002fff10006000e00150023000afff2fffe000a00010000ffd2000dffed0000ffd600070007ffedfffb0035ffe50000000000aefff9fffdfff500000000001cffef00000001ffc5ffebffd00000, 1024'hffa9000e00000000002200000002fffb000cfffbffeffffc000cfffbffee005100140017001fffecfff900000007ffe00000000400010005000e00250023000fffebffee0003fffffffbffe40012fff60000ffcffff70007ffeaffec0038fff00000000000b3ffef0005000a00000000001bfff00000ffe0ffc3ffe5ffd00000, 1024'hffc400090000000000230000ffaa0010000e0006ffb2ffc70030005bfff7003cfff7ffc90048ffed001e00000001ffd3000000030040ffb6ffea0031001a000affa40003ffb6001dffecfffb0003003c0000fff0ffeaffecfff300120019fffa000000000094ffe3ffddffd900000000fff8003c0000ffd4ffbf0027ffc90000, 1024'hffb2000f00000000000d0000005fffe10017ffda00090021ffddffb90018002d00190034ffeffff2ffe20000fff6002e0000fffdffda00500024002c001400240028ffc40054ffe7fff7fff50030ffb10000ffc700020013ffefffd80031000b000000000088ffe9003c002800000000001effb00000ffddffe9ffcfffe50000, 1024'hffa900100000000000160000ffdd001c000a0001ffe5ffcb001fffefffc50047002a00170024ffd5fffb00000015ffc50000fffefffcffe00004001d002c001cffd1ffddffe90016000bffd6001b00020000ffc40000000afff9ffec0035ffd80000000000a3ffcc0003000400000000000f00080000ffe8ffc8fffbffc50000, 1024'hffbc00040000000000140000ffbc0025fffc0002ffe4ffb7001ffffcffbf0040002300160031ffbcfff30000002fffc0000000050002ffcafffe0021002b001cffbbffcdffcc0025fff2ffe6000e00260000ffe8fff40021fff2ffec0030ffc3000000000079ffc1fffc001800000000000000210000ffdaffc8fffdffba0000, 1024'hffdcfffb0000000000200000ffb10022ffe7ffe2ffe4ffc2004a000bffe4002f00100027004dffc7ffd70000000fffc60000000cffd2ffccfffa0032001d003dffbaffc8ffdc0014ffc2ffd2fff9002000000004ffc4001effebffbf002fffc700000000004cffe9ffda000300000000fffa002200000016ffceffbdffca0000, 1024'hffddffef0000000000320000ffb50020ffe3fff10001fff9008bffdf000700320014006f0056fff8ffd20000ffefffbb00000009ffc3ffda00010041fffb0038ffe8ffd3ffde0002fffbffb2fff3001900000011ff89fff9ffd7ff760031ffe80000000000170022ffd2ffe800000000fffe00200000002fffcaff68ffe90000, 1024'hffd4ffe500000000003c0000ffbafffffff7002a000b000e0083ffc8001e003affed008b003d0009ffd20000ffd5ffd300000013000fffe700000049ffde001affe3ffc5ffca0000001effe3fff5002800000025ff80fff1ffc3ff6c0034001300000000ffee0014ffde000f00000000fff500190000ffd1ffb9ff6c00030000, 1024'hffdbffd700000000003d0000ffd5ffe10002002a000c002a004500060008002c000400590036001dfff30000000bfff400000016002600020011003effe0fffcfffaffe9ffc3fffd00240006fff6003b0000004affa70016ffb7ffc0002b000700000000ffef0000fff1001700000000fff100000000ffbeffb1ff9fffff0000, 1024'hffddffd600000000003d0000000affbb001fffe5ffd9001b0010002b000b0020000f003a00380018fffe0000fffb001800000022fff5fffb0024002cffef00170009fff9001cffd200240002002affe50000004affc70007ffbaffe9002d0019000000000006ffd8000f000000000000fff5ffaa0000ffe4ffbeffc100000000, 1024'hffccffe20000000000380000002fffe10040ffe6ff9bfff80009002f0000001f003400230042ffe0001b0000001200290000001c001b000c00210038000c0011000efff1005cffceffecffe8003affa400000023ffcaffdcffd0fff20032fff3000000000028ffda002effef00000000fffdff9f0000fffaffc9ffe8fffc0000, 1024'hffc4fff70000000000280000002f00100033fffdff95ffe500120023ffd7002d0058000e0042ffb800200000003a00070000000a00290013001200280027fffd000ffff3004ffff3fff1ffd00036ffad0000fff4ffdbffeaffe6fff7002fffca000000000055ffda0029ffe2000000000008ffc000000001ffdefff2ffe30000, 1024'hffc1000b00000000001900000022001f0020fffeffb5ffdb0004fffdffc3003d00540010002affab000900000033ffe30000000200140018000800180036000a0009ffe00038000a0001ffd6003affbb0000ffd6fff80003fff9ffef002effc1000000000073ffcb001afffb000000000013ffd60000fff5ffe9fff0ffd50000, 1024'hffbc001500000000001300000017001b000fffffffdaffe8fffbfff3ffca0044003f0009001affc2fffc0000002affde0000fffc0007001f000600180033000e0005ffe0001c000fffffffe0002affd90000ffcc00060016fffefff2002bffc8000000000090ffd7000b000a00000000001bffeb0000ffeaffe5ffecffcb0000, 1024'hffbb00190000000000130000000500070004fff5ffedfff600050002ffdd004500200005001bffe3fff600000010ffd80000fffbfff7000f0004001a002a0015fff8ffef0006000a0000ffe60019fff30000ffc9ffff0018fffcfff30028ffe10000000000a5ffe5fffa000400000000001efff40000ffefffdbffe5ffc90000, 1024'hffb900180000000000150000fffffffe0004fff9ffeffffb00160007ffeb00430011000a001ffff4fff900000002ffdb0000fffcfff9ffff0004001c00220010ffeffffbffff00030001ffe3000efffd0000ffc3fff2000afff7ffee0028fff40000000000aafff4fff9fffa00000000001dfff70000fff2ffd6ffe2ffcf0000, 1024'hffb5001600000000001500000002fffd00050001fff1fffd00180001ffec0042000f0011001ffff5fffa00000004ffe40000fffd000100000006001d00200009ffeafffb0001fffffffbffe4000bfffb0000ffbfffec0003fff7ffea002afff70000000000a9fff5ffffffff00000000001efff80000ffecffd7ffe2ffd20000, 1024'hffb2001600000000001400000009fffd0007fffcfff0ffff0011fffcffee004400150013001cffeffffa00000007ffe50000fffdfffe00030008001d0024000bfff1fff700080001fffcffe3000ffff40000ffbdfff00005fff7ffe9002cfff40000000000acfff30004000200000000001efff00000ffeaffd9ffe3ffd30000, 1024'hffaf00170000000000150000000a00000008fffdffeffffb000efffaffea004700170011001cffebfffa0000000affe60000fffdffff00050009001e0027000bffeffff500090000fffaffe30011fff20000ffbbfff30005fff7ffea002dfff10000000000b3ffef0006000500000000001ffff00000ffe8ffd8ffe5ffd00000, 1024'hffae00160000000000160000fffe00040006fffdfff2fff4000ffff9ffe8004900130010001cffeffff90000000bffe30000fffdfffbfffa0008001f0027000bffe6fff5fffffffefff9ffe1000efffb0000ffbdfff40005fff7ffeb002dfff00000000000b6ffef0004000700000000001dfffa0000ffe7ffd3ffe8ffcd0000, 1024'hffb000160000000000180000fffdffff0009fffbffedfff60011ffffffec004800130011001effe9fffb00000006ffdd00000000fffffff900080021002b0010ffe7fff3ffff0004fff5ffe4000dfffb0000ffbffff20004fff5ffeb002ffff00000000000b4fff10002000600000000001afff50000ffe8ffd1ffeaffd40000, 1024'hffac001800000000001a0000000d0000000afffdffe8fffb0012ffffffe400480021000f0020ffe2fffc0000000cffe10000fffe0002000a000b001e0032000dfff2fff4000e0008fffaffdd0012ffeb0000ffb8fff40007fff4ffec0031ffe90000000000b8ffee0004fffe00000000001dffea0000ffefffd9ffe5ffd90000, 1024'hffa800180000000000190000fff9000f0009ffffffe8ffe30012ffefffce004a002f0012001effd4fff900000016ffd10000fffbfffdfffb0009001d003b0012ffe5ffe3fffd00140009ffda001dfff30000ffb8ffff000efff5ffec0031ffdc0000000000b4ffd800070006000000000015fff90000ffe9ffd6ffefffd20000, 1024'hffb2000b00000000001a0000ffc7001b0003fffdffebffbc0018fff4ffb30041002f001b002cffcdfff40000002cffc600000001fff4ffd4000700270039001fffbbffcfffd20016fffcffe8001e001c0000ffd6fff6001dfff1fff00030ffcd000000000097ffb70008001e000000000004001b0000ffdfffc6fffbffbf0000, 1024'hffcdfff60000000000220000ff9f0020fffbffe1ffdaffa50035ffffffcf00370015002a0045ffcaffe800000012ffbe00000010ffd8ffa7ffff002a00230037ffa1ffc6ffd2000bffe7ffdc0017001d00000003ffd90008ffebffd40031ffd5000000000057ffc3fff6000f00000000fff500290000fffeffc0ffe9ffc40000, 1024'hffe5ffe700000000002e0000ffa400210003fffaffd3ffd5004b000a00010034000c002f004dffdc00010000fffaffbb00000014000dffc2fff5002bffff001cffcbffdfffda000dfff8ffe0000800140000002effc0ffd4ffe3ffbf0022ffe80000000000060006ffe3fff400000000fff8003600000007ffc3ffd6ffe50000, 1024'hfff8ffe400000000002d0000ffdefffe00000036fffb0019003500090004001f000800240026000c00000000ffffffee0000000d002d0005fffe0016ffe4ffe4fff60005ffdbfffe0010fff6ffed001b00000033ffd1fff0ffd8ffd70013ffff00000000ffe20020ffe2ffff00000000fff900120000ffedffcfffc600060000, 1024'hffe9ffeb00000000002400000022ffce0000000800260046fff2ffe3001b001dfff0002afff60027ffef0000ffe7000f00000010fff2003300210002ffe5fff3002300060016ffe10024fffc0000ffe60000002a00040002ffd7fff0001c001d000000000004001b0002000f00000000000cffcf0000ffefffd9ffcb000e0000, 1024'hffc7fff80000000000230000004affcd0015fff800180038ffdaffe1001e002bfff80022ffef001bffed0000ffeb002e0000000dfff3004f00280019fff50007002dfff20041ffd3fffbfffa000bffc500000007000f000cffd9fff7002e000f00000000004d000f0019001e00000000001bffae0000ffe5ffccffd5fffd0000, 1024'hffb000050000000000240000002effe80011fff1fff90022fff8fffc000f004400060009000a0001fffc0000fff8fffd00000004fff9002c001d001e000b00070018fffe0026fff00003ffdb0007ffdb0000ffe80010000affde00000037fffc000000000099000d000cfff600000000001bffc70000fff0ffbfffe5ffe10000, 1024'hffa8000d00000000002300000004fffb00070007fff80002000a0003ffea0054000a0009001afff4fffa0000000effe3000000030006000c0011001f001c0001fff0fffcfffafffeffffffde000100030000ffd500020014ffe4fffc0039ffeb0000000000bbfff90000000300000000001dffef0000ffdfffbaffe7ffcc0000, 1024'hffa5000d0000000000250000fffdfff80007fff5fff9fffe0008fffbffec005800120012001cfff4fff600000004ffd900000005fff000000012001e00230011ffeefff5fffefffe0007ffdb000dfffa0000ffd20004000effe5fff2003bffef0000000000c0fff4ffff000600000000001dffeb0000ffe9ffbbffe3ffce0000, 1024'hff9f000d00000000002900000000fff7000ffffdffeffffd0008ffffffee0059001000120020fff1fffc00000005ffe10000000600040004001200270025000dffe8fff30002fffafffcffe20010fff50000ffd1fffd0003ffe5fff2003cfff10000000000c4fff10004000a00000000001dffec0000ffddffb8ffe9ffcf0000, 1024'hffbe00090000000000280000ffa2001000120008ffaaffbf0030006afff60040fff1ffbc004dffef002400000001ffd300000004004bffb0ffe90036001c0009ff990007ffaf001cffe4fffd000000430000fff2ffeeffe9fff0001e001bfff90000000000a3ffe2ffdaffd500000000fff700420000ffd0ffb40034ffc50000, 1024'hffa9000e00000000001000000066ffd30017ffd6001e0035ffcdffa8002a00370009003fffe40002ffde0000ffe900350000ffffffd6005f002b002f000c00220030ffc2005affdbfff8fffe002fffac0000ffcc0005000bffebffd300340019000000000092fff700420039000000000029ffaf0000ffd4ffdfffc8ffe40000, 1024'hff9d001400000000001d0000fff6fffb000dfffdffedffef0012fffeffe300510014000f0022fff2fffc0000fffdffda0000ffff0004fffc0009002200210013ffd9ffeefffd0003fffeffe20015fff60000ffbefffefffffff3fff30038fff30000000000c8ffe600010005000000000021fffb0000ffe5ffbdfff3ffc40000, 1024'hffaa00080000000000190000ffc30016fff30008fffaffd30021ffebffcf004c001800150028ffd5fff00000001fffc10000ffffffefffca0007001a00270008ffb7ffe1ffc9001afffcffd2fffd00270000ffd3fffe0013ffedffeb0034ffd90000000000acffe5fffe001000000000000900200000ffe6ffbafff3ffb60000, 1024'hffb8ffed0000000000260000ff82001bffd7fff40039ffb90032ffa4ffcd004100050066002affe0ffbf0000001fffc100000010ff9aff9e001b003100200031ff91ffabffa2fffeffdeffceffee004c00000008ffd9001fffd7ffac003dffd1000000000068ffe60003005200000000fff5003d0000fff5ffa3ffb9ffb90000, 1024'hffb7ffcd0000000000500000ff89fff40003ffcc0016ffd00051ffae000f0041fffd00a9004bfff7ffc90000ffe2ffcb0000002cffa5ffa7002a0066ffff0068ffb2ff8dffd0ffdeffeaffe00018001c00000051ff9dffe8ffaeff780051fffc000000000016ffec000c004900000000ffe9000f0000fff5ff7fff90ffe00000, 1024'hffbcffba00000000006b0000ffbfffe40033000effb7fff60063001b00130042001400790071000000090000fffffff8000000310032ffd20020006dffe0001bffdbffd0fff1ffd30008ffea0020000200000076ff7cffcfff97ffa5004d000300000000ffefffee000a000500000000ffe3ffe50000ffcaff79ffa1fff70000, 1024'hffd8ffc100000000005d0000ffebffed00410027ff890000002b005500070041001f00140059ffea003600000015fff70000002c006bffe50011002fffe4ffde00010013000affe70035ffec0022ffe700000078ffcaffcbffaafffb0032fffb00000000ffe9fff40003ffd300000000ffe6ffcb0000ffc8ff9affed00010000, 1024'hffebffd600000000003d0000001a00000031003dffc20002ffd50037ffe70030001affd10011fff0003000000029001a0000001c006000260012fff8fff2ffbc00100029001dffe10012fff80007ffd600000053002dffe5ffd0003e001cffe100000000fffc00010008fff500000000fffeffd20000ffdbffbc002700060000, 1024'hffe3fff400000000002200000040ffe70017fff7fff9001fffb0001bfffd0022000affc8ffebfffd000c00000005001c0000000e000a0055001ffff30007ffef00230013003cffe9ffe8fff50001ffc10000001f0057000fffe8004b0022ffe4000000000042000b00060000000000000012ffc100000009ffcf002600050000, 1024'hffc9000d00000000001b00000039ffe70007ffd9fff7002affe0001b000500300015ffdc0004fff800020000fffcfff40000ffffffec0045001a0008001d000c0027000b00320005fff9ffde0007ffd00000ffeb0032001bffec00280028ffea00000000008d0010fffcffe200000000001bffca00000019ffd9ffffffef0000, 1024'hffb5001c00000000001a0000001ffff30005fff4fff000110008000fffe40043001efffe0018fff3fffa0000000affde0000fff9fff80024000e0017002d000b000b000200140008000bffde0013ffeb0000ffc20004001efff00003002cffeb0000000000b7fff5fffbffee000000000021ffe00000fffaffdaffe1ffd80000, 1024'hffac001b0000000000180000000bfffe0007fff7ffeffff9000efffcffdf004d00180010001bffeffff50000000bffdb0000fffbfff30006000a001e002d0010fff2fff60006ffff000bffdf0019fff50000ffb8fff80014fff4fff00030fff00000000000c4ffe500040000000000000020ffec0000ffe8ffd3ffdfffcb0000, 1024'hffaa00150000000000190000fff600060007fffefff2ffeb0011fff5ffe40050000f0015001dffeefff600000009ffde00000000fff8fff2000800210028000fffddfff1fff8fffbfff9ffe0000f00000000ffbcfff40005fff5ffe80033fff00000000000c0ffea0004000c00000000001dfffc0000ffe2ffcaffe7ffca0000, 1024'hffab001100000000001c0000fff500050007fffdfff1fff20015fffdffee004e000e00120022ffeffffa00000004ffe000000002fffffff60008002300230010ffdffff4fffafffefff1ffe00008fffe0000ffc4fff2fffefff3ffe70033fff00000000000b6fff3fffe000700000000001cfffc0000ffe8ffc9ffe8ffd00000, 1024'hffab001200000000001d0000000100010007fffffff0fffd00160001ffee004e001300110022fff2fffb00000006ffe20000000000020002000900200022000affebfffa0003fffffff8ffdd0009fff70000ffc3fff10002fff1ffe90033fff00000000000b5fff7fffdffff00000000001ffff50000ffebffcdffe2ffd20000, 1024'hffa9001500000000001c00000007fffe0007fffffff000010012fffeffef005000130011001ffff0fff900000007ffe20000ffff00010006000a00210024000afff0fff800050000fffcffde000cfff60000ffc0fff30007fff1ffe90033fff10000000000bdfff7ffff0001000000000020fff00000ffe5ffceffdfffcf0000, 1024'hffa7001700000000001c00000006fffe00070000fff300000010fffdffec00520012000f001dfff1fff900000006ffe00000fffe00000007000a00200027000affeefff900030000fffcffdf000bfff70000ffbcfff60007fff2ffeb0033fff10000000000c5fff6ffff0003000000000022fff10000ffe6ffccffe1ffce0000, 1024'hffa5001600000000001c0000fffc000200060001fff5fff60012fff9ffe700520011000f001cfff1fff800000007ffdd0000fffefffdfffc000a00200028000bffe4fff6fff90001fffeffdd000affff0000ffbbfffa0008fff1ffed0034fff00000000000c7fff10000000500000000001efff80000ffe4ffc8ffe7ffcd0000, 1024'hffa5001600000000001d0000fffc00010007fffffff2fff6000ffffeffe700530010000f001effedfff90000000affdb000000010000fffc000b0022002b000fffe6fff5fffa0002fff8ffe0000bffff0000ffbffffa000afff1ffef0036ffec0000000000c7fff0fffe000700000000001efff50000ffe0ffc8ffe9ffcd0000, 1024'hffa3001800000000001e0000000dfffd0007fffdfff30004000b0000ffed00560012000c001dfff3fff90000000affe50000fffffffc000b000e0021002a000afff7fffe000afffafffaffda000afff20000ffbcfff8000afff0ffed0035ffed0000000000cffffafffe0001000000000025ffe70000ffe7ffccffddffce0000, 1024'hff9e001a00000000001f0000fffffffe00080001fff5fffa0012fff8ffeb00550010000e001cfff3fff800000003ffe00000fffdfffcffff000d0026002d000dffe8fff6fffdfffefffcffda0009fffb0000ffb6fff80005ffefffea0034fff10000000000d6fff800000005000000000020fff20000ffe5ffc5ffe2ffce0000, 1024'hffa100130000000000200000ffd8000e0005000afff7ffd8001cffebffce0051001a0014001effe0fff80000000bffc40000fffffffdffe1000a001e00340010ffc7ffe5ffdc00130007ffda000b00100000ffbf00040006ffedffef0036ffe40000000000bfffe00001000d000000000011000f0000ffe5ffbcfff9ffcd0000, 1024'hffaffffc0000000000220000ffac001a0002fffffffaffb40013ffe2ffaf0046002c00270025ffcafff40000002bffb500000008ffefffbf000e00200036001affaaffc6ffba001e000cffe70018002c0000ffed0006001bffe3fff60038ffcc000000000084ffb3000f002b00000000fff800280000ffdaffb0000bffc70000, 1024'hffd4ffe50000000000300000ff9300190008ffdaffceff9a001d0006ffd0003a001b00260042ffb2fff000000015ffb40000001effeaffa20005002a00280039ff98ffb4ffc90019ffe9fff1002300200000002bfff0000bffd8ffe90039ffcf000000000035ffadffff001f00000000ffe100280000ffeaffaf000bffd40000, 1024'hffefffd700000000003f0000ffb400250008fff8ffc7ffd500390017ffe80031002c00250050ffce000400000019ffc30000001e0002ffd30004002400090018ffdaffe3ffe90008fffaffd2000f00030000004fffd5ffeaffd5ffd6002bffcb00000000fff1fffaffe7fff000000000ffeb001b00000014ffbfffd8fff20000, 1024'hffebffdc00000000003b00000001fff200110016fff70029001200000014003000090030001f001700010000fffb000100000016001a0020000e001affe6fff2001c00030010ffe0001cfff4000affe700000048ffdaffe7ffd0ffd6001f000300000000ffe6001cfff30003000000000007ffea0000ffedffcaffbc000b0000, 1024'hffd6ffe900000000002f00000042ffc000130013001e005affe0fff3002d002fffe70020fff6003ffffa0000ffe5003400000011000b005100250012ffd8ffe0003200190030ffbd00140001fffcffd500000027fffefff4ffcffff80022002700000000002d002e000d001700000000001effb80000ffe0ffc1ffc400080000, 1024'hffb7fff900000000002a00000040ffbc0010fff4001a0043ffe3fff000350035ffdf0011fff6002ffff10000ffd300300000000cffed003e002a001afff1fffb000c00070035ffcaffe9fff0fff5ffd10000fff50011fff6ffd500010035002900000000008900290016000f00000000001fffb90000fff2ffb5ffdffff70000, 1024'hff9d000400000000002a00000010ffe70007fff40008001e0008fff60011004ffff800140015000efffb0000fff5fff600000006fff3001000210025000f0003fff40002000bffebfff2ffd4fff7fff30000ffdb0004fff9ffdbfff8004000040000000000bf0019000afffc00000000001effe40000fff0ffafffe6ffda0000, 1024'hff9a000900000000002c0000fffcfff9000a0005fffa00000010fff7fff3006100060019001ffff8fff700000004ffe1000000080000ffff00150027001a0008ffe8fff7fff9fff50000ffd9000300000000ffd5fffc0006ffddffeb0042fff30000000000c9fffc0001000a00000000001effeb0000ffd9ffadffdeffca0000, 1024'hff99000b00000000002e0000fffffff9000f0002fff2ffff000a0003fff200630009000e0020fff8fffc00000003ffe2000000080007000600130028001e000affe9fff9fffefff6fffaffdc0007fffa0000ffd400010005ffe0fff40043fff00000000000d1fff9fffe0006000000000020ffeb0000ffdaffacffe7ffcb0000, 1024'hffb9000800000000002c0000ff9a000e00120009ffa7ffc20036007afffd0046ffeaffb30053fff500280000fffdffd0000000050054ffacffe7003b00170009ff95000dffa40020ffe3fffdfff8004f0000fff6ffedffebffec0023001efffb0000000000afffe6ffd1ffcd00000000fff600460000ffcbffaa0037ffc20000, 1024'hffa5000a00000000001400000066ffca001bffce0026003affc2ff9a003a003efffe004cffdc0004ffda0000ffde003600000004ffd2005e00300034000900260030ffb8005cffd5fff600060032ffaa0000ffd400070006ffe4ffcd003a0023000000000091fff9004a0048000000000028ffac0000ffc8ffd5ffc9ffe80000, 1024'hff9a001200000000002600000007ffee000ffffffff10007000a0006fff6005b000a000b0020fffefffe0000fff6ffe700000003000b000e000f0024001b0006ffe3fffc0008fff6fff5ffe3000cfff00000ffc2fffdfffaffeafff6003dfffd0000000000d7fffa00000004000000000027fff10000ffe2ffb6ffecffcb0000, 1024'hff9e00080000000000220000ffc70009ffef000b000dffe8001cffdeffe00057000d0015001fffefffed00000010ffcc0000ffffffe2ffcd001000170022fffcffb7ffedffca000c0004ffc8fff400240000ffce00050007ffe6ffe80037ffec0000000000c8fffffffe000f00000000000f00200000ffe9ffb1ffeaffba0000, 1024'hffa4ffe400000000002e0000ff64001bffda000c0069ffb70013ff61ffc80056fffa00780001fff0ffc200000015ffa900000013ff93ff820029001c001e001bff85ffa7ff7efffd0015ffcfffeb005c00000013000c0008ffcbffb3003fffe1000000000069fff00016007700000000fff100500000ffdaff85ffd8ffc00000, 1024'hffabffbc00000000005c0000ff89ffdf0023ffe60030ffc4ffebff9600020051ffe7008b000ffff4ffe00000ffe6ffd00000003effd7ffb5003e004ffffe004effa5ff82ffbbffdd0000001b00250023000000800006ffe5ff9cffca0058000300000000000dffcd0031008c00000000ffe1000d0000ffabff51fffaffea0000, 1024'hffc6ffaf0000000000750000ffe7ffdd004c0002ff9dffeefff600530005004b001200020046ffe8002c00000002fffc0000003e0053000200290035ffe80002ffe7fff20012ffe00006fff80023ffd80000009f0010ffddff96002d0054ffea000000000000ffde000afff300000000ffe1ffc30000ffd1ff62002000060000, 1024'hffe7ffc90000000000590000fff90011002e000fff7bffe8000b0091ffec00400028ffaa0052ffc3003500000021ffe9000000250067001b0004000dfffaffe2fff200210017000fffedffd40000ffdb000000700023fffbffbe004f003effbb000000000015fff2ffdaffa900000000ffeaffde00000008ff9b002efffe0000, 1024'hfff5ffe700000000003600000000002400090006ffbc000a000e0066ffda003c0039ffbb0038ffe100240000002bffc50000000c0030002efffbfff60002ffe8002100300001001f0020ffccfffffff40000003f00260019ffdf00390025ffb90000000000230006ffc9ffab000000000004fff800000021ffcc0004fff40000, 1024'hffe5fffa00000000001f0000002affe6000400050004003affe2001ffff700360011fff20002001f00010000000dfffb000000060002003b000dfff9fff9ffeb003500250010fff00036fff5000bfff00000001400190027ffe70018001afffa0000000000440004ffecfff4000000000019ffce0000ffebffdeffdbfff40000, 1024'hffca000500000000001800000039ffc90007ffec001b0036ffd7fff300250030ffe50007ffee0024ffec0000ffe0002400000007ffdd002e001e000c000200010014000b002dffd3fff5fff7fffbffda0000ffe80013000affe800000024001e0000000000800016000d001500000000001effba0000fff1ffd4ffdffff70000, 1024'hffa9001000000000001f00000029ffe0000cffeb000d0027fffcfff1001f003ffff4001200060015fffb0000ffe9000a00000002ffed001f0020002500190009000600050024ffe1ffe4ffdffff9ffe10000ffc6fffffff1ffe7fff40032000f0000000000b9002300120002000000000023ffd70000fffbffc9ffe5ffef0000, 1024'hff9c001700000000002200000010fff3000c0004fff600080013fffafff50051000b0011001afffefffc0000fffdfff00000fffe0006000c0012002500270002ffebfffe000afff6fff9ffdc0007fff10000ffb3fff4fffcffeaffee0037fffe0000000000d3fffe0008ffff000000000022ffec0000ffe5ffc7ffe4ffda0000, 1024'hff9c001600000000001f0000fff5000500070001fff3ffed0010fff6ffdc005800160011001fffeafff90000000effd60000fffffffffff6000c00210030000bffd9fff1fff50004fffeffdc000f00000000ffb8fffe0008fff0fff10039ffea0000000000d4ffe70004000a00000000001effff0000ffdfffc3ffefffc80000, 1024'hffa200120000000000200000fff300060009fffaffeeffe9000afffbffdd0059001800100022ffe5fff90000000fffd400000003fffbfff6000b0021002d0013ffdcffedfff80003fffaffe00014fffd0000ffc500000009fff0fff1003affe60000000000caffe40002000d00000000001efffb0000ffe1ffc0ffefffc30000, 1024'hffa300100000000000220000fffe0002000afffaffedfff6000cffffffe60058001700100023ffebfffa0000000bffdc00000003fffb0000000d00220027000fffe8fff50003fffcfff9ffda000ffff40000ffc8fffb0006ffeeffee003affe80000000000c6ffef00000006000000000020ffef0000ffe8ffc0ffe5ffc90000, 1024'hffa0001100000000002300000003fffd000bfffbffeffffe000effffffef0059001200120022fff0fffb00000008ffe000000002ffff0003000e00260026000cffebfff70004fffbfff9ffdc000cfff60000ffc5fff60004ffebffec003affef0000000000ccfff600030005000000000021ffee0000ffe4ffbfffe2ffcb0000, 1024'hff9e001300000000002400000002fffa000afffffff0ffff000f0000ffee005b000f00100022fff4fffb00000005ffe10000000200010002000e002400270008ffe7fffb0002fff9fffaffdc000bfff70000ffc0fff60001ffebffed003afff30000000000d4fff800010004000000000023fff00000ffe3ffbfffe2ffcc0000, 1024'hff9c00130000000000240000fffcfffd00090000fff3fffa0010fffbffea005a001100100021fff2fffa00000004ffde00000001ffffffff000e00240029000affe0fff7fffdfffcfff9ffdb000afff90000ffbefffa0000ffecffed003afff10000000000d5fff500010007000000000021fff50000ffe5ffbdffe6ffcc0000, 1024'hff9b00130000000000240000fffbffff0008fffffff4fff8000ffffcffe9005c000d00110021fff3fff900000008ffdc00000002fffffffd000e00250029000cffe0fff7fffbfffbfff7ffdc000afffd0000ffc0fffb0004ffecffef003cffef0000000000d7fff400000008000000000022fff70000ffe0ffbcffe7ffc80000, 1024'hff9c001200000000002400000000fffd0007fffffff80002000bfffcfff1006000080010001efffafff900000007ffe000000002fffb0000000f002400240007ffeafffffffdfff4fffbffd90005fffd0000ffc3fffa0004ffebffed003bfff20000000000dafffeffff0007000000000025fff00000ffe0ffbaffdfffc80000, 1024'hff9a00120000000000260000fffbfff700080002fffd0001000efffafff8005e00000010001c0000fff80000fffbffe600000003fffdfffd0010002700220008ffe0fffdfff8fff2fff4ffddffff00010000ffc0fff9fffdffe8ffeb003bfffb0000000000dd0002ffff000b000000000023fff30000ffe0ffb5ffe2ffce0000, 1024'hff9700110000000000280000ffeffffa00080002fff9fff60016fff8ffe9005a000d00120021fff4fffa0000fffcffd800000003fffffff700110024002a000cffd4fff4fff20001fff9ffd9000400000000ffbffffefffcffe7ffef003efff30000000000d7fff6ffff000700000000001dfffc0000ffe8ffb4ffedffd20000, 1024'hff9c000a0000000000280000ffd40010000a0005ffedffd20016ffe5ffc40057003000190020ffc6fffa00000013ffb300000004ffffffe0000f001b003d0013ffc7ffd5ffdc00260014ffd5001600080000ffcd0013000dffe3fff40041ffd50000000000b5ffd00007000f00000000000600080000ffe2ffb30004ffd30000, 1024'hffb0fff700000000002c0000ffaa002f00090003ffe0ff980012ffeaff93004a0048001e002dffa0fff400000044ffa60000000efffbffc3000e002400480028ffa8ffb0ffb700350008ffe3002500290000fffc00180033ffdc00000044ffa900000000007bff94000c002a00000000ffe8001f0000ffd0ffac0018ffc60000, 1024'hffd1ffe00000000000360000ff9500340007ffd9ffccff9100130001ffac0049003600240042ffa6fff100000036ffa10000001fffddffad000a00200031003cffb6ffb7ffcd001c000cffda003000150000003e00040023ffd7fff10040ffa900000000002eff9bfff9001600000000ffe4001b0000ffefffae0002ffcd0000, 1024'hffeaffd40000000000430000ffc2001b001bfff3ffc6ffd70015001afff00041002500210040ffd3000900000016ffca000000230011ffe2000500290004001bfff2ffdffff3fffd000bffea001efffc00000061ffe6fff3ffccffe3002dffce00000000fff0ffebfff0000600000000fff000040000fff4ffafffe3fff20000, 1024'hffebffdc0000000000420000001bffd8001d001affef0045ffef002100210037000100060014002700180000fff5000e00000019003000330016000bffe2ffd200290029001cffd40025fffd0006ffde0000004efffbffdcffc80006001b0014000000000003002ffff8fff600000000000dffd80000ffebffbfffdd00130000, 1024'hffcfffed00000000003100000050ffb400120011002b0059ffc5ffeb0025002dffe8000affe30042fff70000ffde004400000010fffa005b00300000ffe6ffd4001d001f003dffb6fffffffcfff5ffc4000000120023fff2ffd100140027002b000000000053002f0018001e000000000020ffb40000fff2ffbeffe1000f0000, 1024'hffa3fffb00000000002c00000030ffc3000effda00240036ffd3ffd900320041ffe30017fff00025fff00000ffd8001c0000000dffd5002c0034001d0005000afffefff5002fffd2ffe7ffe80000ffd10000ffef0027fff3ffd60008004000210000000000ab00220023001900000000001effcb0000fff2ffacfff6ffee0000, 1024'hff95000100000000003200000002ffee000efffb0001000c0000fff70001005fffff0013001a0003fffe0000fffeffeb0000000bfffc0008001f002700150005ffe7fffb0002ffecfff4ffdafffffff70000ffe2000bfff8ffd8fffb0046fffa0000000000cd000b000b000b000000000020ffea0000ffe3ff9fffeeffcd0000, 1024'hff93000500000000003300000001fff300120000fff0000100050008fff300670006000c0023fffdffff00000003ffe60000000b000700060017002800190007ffe5fffe0001ffeefffaffdb0007fff70000ffdb00060001ffdbfffc0048fff30000000000d9fff900020006000000000022ffe50000ffdaffa0ffebffc70000, 1024'hffb500040000000000300000ff97000c00170005ff9bffbe0034008600020049ffe7ffab005afff2002e0000fffbffd200000008005bffa8ffe7003f0015000aff8d000effa5001effdafffefff9004d0000fffcffefffe3ffea002a0022fffc0000000000b7ffe5ffd2ffc900000000fff500450000ffcaffa00041ffbe0000, 1024'hffa0000700000000001700000067ffc80020ffcb00270034ffb8ff8e0039004000000055ffd6fff9ffd60000ffe1003600000008ffd1005e0035003a000f002e002dffa7005cffd8fff2000c0038ffa90000ffd9000e000dffdfffcd0041001f000000000091ffee00540058000000000022ffa60000ffbaffceffcfffea0000, 1024'hff96000f00000000002c0000000ffff30011fffcffed000800040009fff20063001000090021fff9ffff00000002ffe700000006000700130014002500210007ffeeffff000efff3fff6ffdb000dffeb0000ffc800030002ffe5fffa0044fff20000000000e0fff900010001000000000027ffe40000ffe1ffb2ffe9ffcb0000, 1024'hff9700040000000000280000ffc1000fffef000d0016ffe50017ffd3ffe4006300030017001afff9ffea0000000effd100000001ffdbffc800130019001efff9ffb7fff0ffc6fffe000affc1ffef00260000ffd400090003ffe1ffe3003affed0000000000d00004fffe001500000000001100200000ffe4ffa6ffe4ffba0000, 1024'hffa1ffe00000000000360000ff50001fffdf001a0072ffae000fff54ffcf0060ffeb0072fff4fff2ffc60000ffffff9a00000018ffa2ff790027001500180017ff78ffa5ff6c0003001effd2ffe200640000001c0025fff6ffc5ffb90042ffe8000000000063fffb000f007d00000000ffed005f0000ffd3ff72ffeeffcc0000, 1024'hffafffbf0000000000610000ff98ffe00027fffa002cffd2ffd7ffad00020058ffdf0060ffffffe8ffed0000ffdcffc10000003f0009ffdf0037003bfffe003cffaeff8fffbbfffa000000280019001e000000870036ffebff9dfff5005bfffa00000000000bffd4001d007e00000000ffe400130000ffa2ff4e0023fffc0000, 1024'hffcdffbe00000000006e0000001bffd90045fffbff990012ffd90083fff00050002cffc7003bffe2003400000012fff0000000320061004d00230019fff4fff50014000f002700010015fff90023ffc90000008f00410011ffa000670055ffd1000000000024ffd7fff4ffd000000000fff2ffaf0000ffe3ff74003100070000, 1024'hffd6ffd800000000004b0000001cffff0022ffe7ff89fff7fff80090ffbf0042005cffb20052ffc5002500000042ffe40000001800240031001200060016fff6000a001d00270015000effc80020ffd000000047002c003affc5005c0047ffab00000000005cffc3ffebffab00000000fff7ffb80000001affaa0015ffe30000, 1024'hffd2ffee0000000000340000ffee00220014ffc8ff97ffc9001f0046ffca00460050fff50057ffac000800000027ffba00000013fff2fff300020019002a002ffff0ffe9001c001b0005ffc20035ffd400000018fffd001affe200040041ffb400000000005dffbbffedffc700000000fffcffe00000001fffc8fff2ffd40000, 1024'hffd2fff700000000002c0000fffa003100140006ffb9ffe9002a0018ffd9005000410014003fffc6000a00000027ffc50000000a001e0009fff8001c00160007000dfff7000f000d0017ffcb0020ffe300000004ffe20002ffebffdc0032ffc300000000004affe8ffedffe100000000000dfff30000fff8ffd4ffd0ffdf0000, 1024'hffc9fffe00000000002100000024fffe0007001700060022ffffffe9ffed004900220025000afff8fff100000014fff60000000500050036000d0010000afff2001bfffb0011fff60017ffe60008ffea0000ffecfff6001bffe7ffe00030ffea000000000067fffc0002001500000000001cffd80000ffdfffd4ffbfffec0000, 1024'hffab000800000000002300000035ffd6000dffe1000d002dffe8ffe70019004d0001002300010008ffea0000ffe9000600000009ffe60033001e0020001600170012ffed002cffeb0000fff10014ffd40000ffd700060010ffe2ffe9003d000e0000000000a8fffb00110018000000000022ffc00000ffdeffcbffd3ffee0000, 1024'hff9800110000000000290000001cfff1000dfff9fff3001300060000fffe005b000f000b001cfffffffb0000fffefff700000002ffff001b0016002600230006fff900000018fff0fff7ffd7000affe30000ffc0fffd0000ffe6fff0003efff90000000000da00020004fffd000000000026ffdc0000ffe7ffc1ffddffd80000, 1024'hff9300170000000000260000fff6fffe00060003fff7fffa0012fffaffe70061000f000d0021fff5fff900000004ffd90000fffffffffffc000f0025002d0008ffddfff9fff6fffefffcffd60007fffe0000ffb8fffd0002ffebffee003cffef0000000000e7fff7fffc0005000000000023fffa0000ffe2ffb9ffe6ffc80000, 1024'hff9700150000000000260000ffeffffe00080000fff7fff2000ffffaffe20061000e00110021ffeefff900000006ffce000000020000fff7000e0025002e000effd8fff2fff00003fffdffdf000b00050000ffc000000006ffe9fff2003dffed0000000000dfffefffff000d000000000021ffff0000ffdeffb4ffedffc40000, 1024'hff9a00110000000000280000fffcfff9000bfffdfff2fffa0007fffeffe400610013000f0020fff0fffb00000009ffd600000004fffe000000110021002b0009ffe2fff7fffcfffd0001ffdd0010fffa0000ffc600030007ffe7fff7003fffee0000000000dbfff000030009000000000022fff30000ffe0ffb5ffebffc70000, 1024'hff9900100000000000290000fffffff9000cfffbfff0fffa0005fffdffea00610012000d0020ffeefffa00000005ffdd00000005fffd000200120023002a000bffe1fff50001fffafff9ffdc000ffff40000ffc600040003ffe7fff40040ffef0000000000dcfff10003000a000000000021ffee0000ffe1ffb5ffebffc90000, 1024'hff97001100000000002a0000fffdfffd000bfffdfff2fffc0009ffffffeb00630010000c0021fff2fffc00000007ffdb00000004ffff000100120025002a0009ffe3fffafffefff9fff8ffd8000afff80000ffc500020002ffe7fff40040ffed0000000000e0fff700000006000000000022fff20000ffe2ffb4ffeaffc90000, 1024'hff96001200000000002a0000fffbfff9000afffffff5fffd000afffdffeb0064000e000e0020fff4fffa00000004ffdb00000004fffe000000120024002a0008ffe1fff9fffcfffafffbffd90009fffa0000ffc300000003ffe6fff20040fff00000000000e3fff800000008000000000023fff30000ffe1ffb3ffe7ffc90000, 1024'hff94001100000000002b0000fff8fff8000afffdfff7fffc000afffcffec0064000d00100021fff6fffa00000003ffda00000004fffefffe00120026002a000affddfff7fffafffafffaffdc000afffc0000ffc400000001ffe5fff20040fff20000000000e3fff70001000b000000000023fff70000ffe0ffb1ffe9ffc80000, 1024'hff96000f00000000002c0000fff7fff8000bfffefff5fffc0009fffcffec0065000c00100020fff5fffb00000003ffd700000005fffefffb0012002400290007ffdcfff9fff8fff9fffdffdb000afffd0000ffc700020000ffe4fff40041fff30000000000e1fff70002000a000000000021fff60000ffdfffaeffebffc90000, 1024'hff96000d00000000002d0000fff9fff7000cfffffff6fffd0005fffcffed0065000b000f001ffff5fffc00000004ffdc000000070000fffe0014002400280006ffdcfff9fff9fff7fffaffdd0009fffc0000ffca0004ffffffe3fff60042fff30000000000e0fff70004000d000000000021fff40000ffddffadffedffcb0000, 1024'hff93000e00000000002e0000fffdfff3000dfffcfff500000001fffeffee0065000e000c001ffff7fffd00000002ffe000000007ffff000200160023002a0007ffe0fffa0000fff6fffaffdc000cfff40000ffc90007fffdffe3fff80042fff30000000000e3fff80003000b000000000023ffef0000ffe0ffafffeeffcd0000, 1024'hff91001000000000002e0000fff2fff9000d0001ffeffff30007fff9ffe00060001b000a0021ffe5fffd00000007ffd4000000050000fffa001600240035000cffd8ffeefff70006fffdffd7000efff70000ffc7000d0001ffe3fff90041ffe70000000000e1fff00003000b00000000001afff20000ffe3ffaefff5ffcd0000, 1024'hff94000900000000002e0000ffcf0018000b0009ffedffc20013ffe6ffb00059003400130025ffc7fff900000020ffb700000005fff9ffe1001400200041001bffbfffd2ffda001d000cffd1001900080000ffd3001c0011ffe2fffc0044ffc80000000000c3ffc80007001400000000000900080000ffe5ffa80006ffc30000, 1024'hffa8fff300000000002e0000ff9c0033000bfffdffe4ff900010ffe3ff940054003b0023002bffaafff40000003eff9c0000000ffff1ffb4000f00240040002bffa8ffb3ffb300290014ffda0025002a00000006001d002cffda00000048ffa900000000007eff96000b002900000000ffec00200000ffd1ff9a0019ffbd0000, 1024'hffd3ffde00000000003a0000ff96002d0010ffe5ffc1ff9700110012ffbc004d002a00180042ff9afffb0000002fff9c00000024fffeffb200070027002c0035ffb7ffb9ffc400260001ffe7002300220000004800080020ffcefffc0042ffab00000000002fffa8fff7001800000000ffdf00170000ffdfff9e0010ffd30000, 1024'hfff1ffdb0000000000480000ffe5001c001efffaffb4ffec00140040fff20044002bfff9003effd1001600000015ffc900000020002900050001001a000b000b000affff00040009000dffe20015ffee00000055fffcfffcffcc0001002fffca000000000002fff6ffdfffde00000000fff3fff100000001ffbbfff000050000, 1024'hffdeffe900000000003a00000043ffeb0010001d0008004affebfffefff80041002200100001001d000100000009000e0000000f000c0060001efff9fff4ffd3004300250034ffd80031ffdb0006ffc40000002100100008ffd20001002cfff400000000002c001dfffafff600000000001cffbe0000ffffffd0ffc100150000, 1024'hffadfff700000000002d00000043ffc20010ffeb00300040ffc3ffc500240048fff40029ffe10024ffe10000ffdf00270000000effdc004d00300017fffe00050018ffe70035ffd20009fffa0011ffc80000fffa00260010ffd2fff7003e001d00000000008600060022003500000000001fffb80000ffd4ffb8ffd9fff90000, 1024'hff97fffe00000000003500000010ffdb0011ffe7000b001affe7ffef000f005ffffb0013000b0008fff80000ffebffef0000000fffee001a002600210013000effeffff20012ffebfff9ffe5000affe50000ffec0020fffcffd40004004a00060000000000c7000600100014000000000020ffdd0000ffe4ff9dfff6ffd80000, 1024'hff90000300000000003800000006ffeb0012fffcfff1000cfffa000afff6006c000a00050021fffb000200000001ffe30000000c00090011001b0022001bffffffe600000007fff3fffdffdb0009ffef0000ffe00012ffffffd70007004bfff40000000000e0fffe00040004000000000024ffe70000ffdeff9cfff3ffc90000, 1024'hffb400040000000000350000ff93000600180001ff96ffbe002e00900002004cffe9ffa1005dfff000300000fff8ffcd00000009005fffaaffe6003f0019000bff84000cffa20024ffd70005fffe004e00000000fff7ffe3ffe800340023fffe0000000000c0ffe2ffcfffc900000000fff4004c0000ffc9ff9b004bffbb0000, 1024'hff99000700000000001900000069ffc50020ffca002e0035ffb0ff81003800430001005cffd1fff4ffd10000ffe3003700000009ffce0064003a003e00140032002dff9b005dffdafff0000f003bffa70000ffda00130012ffdcffcb0045001c000000000097ffeb005a0065000000000022ffa40000ffb2ffcaffceffe90000, 1024'hff90000e0000000000310000000cfff20010fff9fff1000900000006fff1006a000e000a0021fffbfffd00000003ffe20000000700010013001700270024000affeffffe000cfff1fffaffd9000effec0000ffcd00080004ffe1fffb0047fff00000000000eafffb00000004000000000029ffe30000ffe0ffaaffe6ffc70000, 1024'hff94ffff00000000002e0000ffb80010fff300100019ffde0017ffceffdf00680002001b0018fffaffea0000000bffcb00000003ffdaffc30015001b001dfff9ffafffedffbcfffb000fffc1ffee002c0000ffda000e0002ffdaffe5003fffed0000000000d1fffe0001001b00000000000d00210000ffe2ff96ffe8ffbc0000, 1024'hff9effda00000000003d0000ff56001bffee0013005dffa7000aff69ffc80063fff4006dfffcffe8ffd200000002ff960000001fffb4ff7e00290019001a001dff76ffa3ff7200070020ffdbfff0005d00000025002bfff7ffbfffcb004cffe5000000000064ffe40016007800000000ffe900550000ffcbff680002ffd00000, 1024'hffadffc00000000000620000ffbaffdf0034fff00001ffd5ffccffddfff8005cfff900440011ffdcfffe0000fff3ffd100000040001dfff30034003800050036ffc1ffa1ffdefff9fffb0025002c0001000000820036fff4ffa2000d0060ffec00000000001fffc1001e006300000000ffebfff70000ffa3ff5b002dfff50000, 1024'hffc5ffce0000000000650000003fffe00042fff0ff86001bffd8008cffee00570041ffba0044ffd500320000001cfffc0000002a00520060002100150001fff5002d001c0051fffa0007ffe00029ffa40000006b003a0013ffb0005d0055ffc3000000000051ffe0fff0ffbc000000000004ff920000fffaff8c001bfff90000, 1024'hffb8fff2000000000042000000330003001efff1ffa3000dfff4005bffc300560064ffc4003effc7001f0000003cffdb0000000a00160042001900060026fff10028001b003700140023ffb50024ffbc000000140031002cffd000400045ffaf00000000009affe1fff4ffb400000000000fffb000000018ffb5fffdffd70000, 1024'hffaa000400000000002f0000ffe8000e0011ffe7ffc6ffca00060018ffb2005300460003003affbafffb0000002fffc200000009fff5fff800100025003f0026ffdbffd4fffd00190006ffd90033fff00000fff0000c002bffe100080042ffbb0000000000aaffb100020001000000000008ffed0000ffeeffb6fff9ffbc0000, 1024'hffb600020000000000300000ffd8001c0013ffe3ffb5ffbf0028001fffbf0051003f0014004dffb5fffd00000022ffb20000000dfff8ffe20005002e00380032ffd8ffd6fffe0015fffbffd0002ffff10000fff3ffeb0014ffe4ffec0041ffbd000000000090ffbffff6fff2000000000006fff60000fffeffb9ffe8ffc20000, 1024'hffb4000100000000002f0000000d001600150000ffcefff50021fffaffcb0059004b00300037ffc7fffe00000029ffc60000000900010012000f00220029000e0011ffea001c0005001dffc5002affd70000ffe9ffe4000effe0ffd70041ffc7000000000084ffe20005fff6000000000017ffd70000fff6ffc7ffc1ffd40000, 1024'hffa0000800000000002d00000031fff2001cffffffe70011fff5ffe8ffed0060002a002e0018ffe0fff300000014fff700000009000900340019002d0024000b0014ffdf002dfff1000cffe8002cffcd0000ffdafff20014ffdeffdd0044ffe90000000000adffe00019001d000000000022ffc20000ffc7ffc3ffc7ffd60000, 1024'hff96000e00000000002e00000017fff50011fff8ffee0009fffbfffefff300670014000c001dfff7fff900000007ffef00000005fffb00180016002700250008fff7fffa0016ffecfffeffd90014ffe30000ffcb00030007ffe3fff20042fff10000000000e1fff600070008000000000027ffda0000ffdeffb5ffdcffca0000, 1024'hff90001100000000002d0000fff4fff9000a0002fffafffd000bfffcfff100680004000c001f0001fffb0000ffffffdf00000004fffcfff80013002800260006ffdafffffff4fff0fff7ffd6000200010000ffc20001fffbffe5fff20041fff60000000000f00001fffe0009000000000024fff70000ffdfffa9ffe8ffc70000, 1024'hff90001100000000002d0000fff1fff4000a0003fffbfffd000dfffefff100660002000e0020fffbfffc0000fffcffda000000060003fff70014002700280007ffd6fffcfff1fff8fff5ffdc000000040000ffc30001fffbffe2fff40042fff70000000000ebfffefffe000b000000000022fff80000ffddffa9ffeeffcb0000, 1024'hff91001100000000002e0000fffbfff7000b0001fff6ffff0008ffffffed0067000b000a001ffff6fffd00000004ffda000000050003ffff00150024002b0004ffe0fffdfffafffafffcffd80006fffc0000ffc500070001ffe1fff90042fff10000000000e9fffc00000006000000000022fff30000ffdeffaeffeeffcb0000, 1024'hff92001100000000002e0000fffafff9000a0001fff9fffc0004fffaffe70068000d000c001dfff4fff900000007ffd900000005fffd000200150024002d0007ffdefff8fff9fff9fffaffd90008fffc0000ffc600090006ffe3fff80043ffed0000000000ebfff80001000d000000000023fff40000ffdeffacffebffc70000, 1024'hff90001000000000002f0000fff8fff7000bfffbfff8fffc0006fffcffec0069000a000e001ffff7fff900000002ffd800000006fffaffff00150027002c000dffdefff7fff9fff8fffaffd90009fffc0000ffc700070004ffe2fff60045fff00000000000edfff80000000b000000000023fff20000ffdfffa9ffeaffc80000, 1024'hff8f000f0000000000300000fff8fff8000b0000fff7fffe0009fffeffec006b000a000e0021fff8fffb00000004ffd900000006fffffffe00150027002a0007ffdffffcfff7fff6fffcffd70006fffe0000ffc700040002ffe0fff50045fff00000000000edfffaffff0009000000000023fff10000ffddffa8ffe8ffc90000, 1024'hff8f000f0000000000310000fff6fff5000c0000fff7fffe0006fffeffee006b0008000c0020fff8fffc00000001ffda000000070001fffd00160027002a0006ffdcfffbfff6fff6fffcffda0007fffe0000ffc90006ffffffdffff70044fff30000000000edfffa0000000b000000000022fff30000ffdbffa7ffecffca0000, 1024'hff90000f0000000000320000fff4fff6000c0002fff7fffb0006fffeffea0069000b000a001ffff6fffc00000002ffd8000000070001fffc00160025002d0006ffd9fffafff5fff9fffaffd90006fffe0000ffc9000a0000ffdffffa0044fff00000000000ebfffaffff000b000000000020fff50000ffdeffa7fff0ffcc0000, 1024'hff90000f0000000000320000fff7fff7000cfffffff7fffc0003fffdffe9006a000c000a001efff4fffc00000004ffd6000000070000000000170024002e0007ffddfff9fff8fffafffcffd90009fffb0000ffcb000d0002ffdffffc0045ffee0000000000eafff80000000a000000000021fff40000ffdeffa8fff1ffcb0000, 1024'hff91000f0000000000320000fffcfff8000d0000fff7ffff0000ffffffeb006d000a0008001cfff7fffc00000005ffd8000000070001000400160024002b0005ffe3fffdfffafff6fffeffd90008fffb0000ffcc000e0005ffdffffd0045ffee0000000000ecfffaffff000a000000000023fff00000ffdbffa7ffeeffca0000, 1024'hff90000f0000000000320000fffcfff0000dfffefffa0007fffc0001fff1006d00060006001afffbfffe00000000ffd9000000070001000500170023002c0002ffe20000fff9fff7ffffffdc0005fffc0000ffcb000e0002ffdf00000044fff40000000000f2ffff0001000b000000000024fff00000ffdcffa5fff0ffce0000, 1024'hff8c000c0000000000330000fff1fff6000c0000fffdfff10002fff2ffdd00690014000b001dfff4fffa0000fffdffd600000007fff900000018001c002d0009ffcdfff2fff7fffc0002ffd9000efff50000ffc60018fffbffdffffe0047fff10000000000ecffee00050010000000000023fffa0000ffe9ffa3fff8ffca0000, 1024'hff8d00010000000000320000ffbe000e000c0000ffefffc4000affe3ffba005f002e00160024ffc9fffa00000015ffaf00000009fff9ffd500150021003c001affacffcaffce0021000dffd6001b000e0000ffdd0024000affdf0002004bffd00000000000c7ffc5000a001d00000000000400150000ffdcff970015ffc40000, 1024'hffacffef0000000000350000ff9a0024000bfff5ffd5ff9d000cffffffa10055003c00160038ff98fffc0000003dff92000000150000ffb6000e0025004a002affa1ffb5ffb2003c0003ffe60020002d00000012001c002affd4000b004affa9000000000082ff9d0006002500000000ffe7001f0000ffd3ff970024ffc30000, 1024'hffd1ffe50000000000420000ffcd002f001dffdbff9fffa0001d0032ffab004a004f000d0054ff91000000000036ffaa000000210001ffe50008002b003b0042ffd5ffc4fff90021fff5ffd80036fff10000003000010029ffd10001004dff9c000000000046ff9afff4fff600000000ffeaffeb0000ffffffaefffeffdd0000, 1024'hffc8ffe900000000004000000024002c001cffefffbafff70019000affc6005c0063002a003dffc3000000000036ffcf00000014fff9003200120018001d0013003afff20040fff9002dffae0037ffb000000019fff1001affd6ffdd004cffab000000000045ffd8fff9ffdb000000000011ffba0000000effccffb3ffef0000, 1024'hffa7fff400000000003600000035ffff001d0007fff60018fff0ffceffec0067003a0041000fffe4ffeb00000019fffd0000000e00000047001d0029000d0008002bffd5002fffeb0026ffde002dffc50000fffcfffa001effd2ffcd004bffde00000000007dffdf0019002800000000001dffb70000ffc5ffb8ffb0ffdf0000, 1024'hff93fffe00000000003900000014ffe40016fff4fffd0011ffeaffedfffd006d000e001f0012fff7fff10000fffaffee00000011fffb00220020002700170011fff8ffe40014fff00008ffe8001affe00000ffed0013000fffd2fff20050fff70000000000c4ffeb000c001f000000000020ffd00000ffcaffa0ffe0ffd20000, 1024'hff8d000400000000003b00000006ffef0011fff9fff1000cfff90009fff60073000f00040021fff7ffff00000003ffdf0000000c00030012001c0024001f0003ffedfffe0007fff5ffffffd50009ffee0000ffe100150006ffd40003004effed0000000000e7fffeffff0003000000000023ffe10000ffdeff9affedffc80000, 1024'hffb1000600000000003a0000ff8c0006001a0004ff93ffbc0034009800020050ffe5ff9e0061fff200320000fff6ffc90000000a0066ffa7ffe60046001b000dff81000dff9a0025ffd70006fffc005600000002fff3ffe4ffe400350024fffe0000000000c8ffe2ffcaffc600000000fff200500000ffc4ff95004bffbb0000, 1024'hff93000600000000001b0000006effbf0023ffc60034003bffa6ff77003d004800000063ffcbfff5ffd00000ffe200390000000affcb0068003f0041001600320031ff960060ffd7fff40013003fffa40000ffdb00160012ffd8ffca0048002000000000009effea0063006f000000000023ff9f0000ffaaffc5ffceffea0000, 1024'hff8c000b00000000003600000007ffed0013fff9fff30007fff70004fff3007000090008001efffeffff00000000ffe30000000a0002000d001a002600250005ffe6ffff0008ffecfffcffdd000fffee0000ffd1000ffffeffdc00010049fff60000000000f2fffa0005000b000000000028ffe60000ffdaffa1ffefffc80000, 1024'hff90fffc0000000000340000ffba000afffd000e0012ffdb000bffd0ffd70069000e00170016fff1fff20000000affc600000007ffe0ffc7001a00180026fffaffabffe9ffc100000011ffc5fff700210000ffdd001dfffcffd7fff30044ffea0000000000d5fff50009001f00000000000a001b0000ffe4ff8efffbffc40000, 1024'hff96ffdf0000000000400000ff7800150004000a0036ffa6fff3ff8bffb90066001000510002ffd2ffe80000000eff9800000020ffd4ff9b002a0015002b001eff88ffa7ff9400130025ffe6000f00390000001f0041fff8ffc2ffee0051ffda000000000076ffc7001f006700000000ffee003b0000ffc5ff700024ffd10000, 1024'hffabffce0000000000580000ffdffff3003cfff0ffdaffcbffb70001ffd60063001a00140015ffc2000e00000015ffd100000036002e000c002b002700170027ffd6ffb8fffd000000000018003dffe40000006800510007ffb50033005dffcd000000000047ffa9001d004700000000fff7ffe20000ffaaff6f0044ffe20000, 1024'hffbeffde0000000000520000004dfff20036ffe7ff980016ffc40078ffdd00610048ffb30035ffd4002900000033fffa0000001f002e00610020000a000efff4003600230056fff20003ffd10027ffa500000046004a0026ffc500600053ffb4000000000088ffe2fff8ffc6000000000016ff9200000002ff980016ffdc0000, 1024'hffa6fffe00000000003900000038fffe001affe3ffc10014ffeb0038ffe400670040ffd6002bffde00100000001fffe400000008fff90039001a000e0022ffff00240018003bfffc0013ffb6001affbd0000fff2002e001dffda0026004affca0000000000d0fff6fffbffcb000000000021ffae0000000fffafffefffcd0000, 1024'hff91000b00000000002f0000ffec000a000efffeffe9ffe40006fffdffd00069002500080025ffdcfffd00000019ffcb00000005fffefff8001300250034000effd9ffeaffef00090006ffd20013ffff0000ffd000110012ffe1fffe0047ffd60000000000e1ffdd0004000a000000000018fff60000ffdeffa6fff6ffc10000, 1024'hff9800070000000000310000ffd80007000ffff4ffe0ffd1000f0009ffc60061002700120033ffd2fffb0000001affc00000000cfffcffe50011002b003a0021ffc6ffddffe6000ffffaffde001b00080000ffdb00050015ffdffffc0049ffd20000000000ceffc900010011000000000010fffd0000ffdfffa5fffbffc10000, 1024'hff9b00050000000000340000000200060017ffebffd0ffea00090007ffd10066003700190034ffcd00000000001dffc70000000dfff90001001600240037001afff4ffea00160003000cffcd002affdb0000ffdf0001000cffdefff3004bffd00000000000c1ffd70007fffd00000000001affd80000ffedffb4ffe5ffca0000, 1024'hff94000a0000000000330000001c0004001d0000ffd9fffbfff9fffaffdd006d003000150024ffd800000000001fffe400000008000c001e0017002b003000070002ffed001ffff40005ffd60025ffd60000ffd40002000affdffff00048ffd80000000000d3ffe40011000d000000000023ffd10000ffd5ffb3ffdeffc80000, 1024'hff90000e00000000003100000003fffd00110000fff0fffafffafffbffe4006f00140008001dfff1fffc0000000cffe000000006ffff000a00160025002b0004ffe6fff90003fff00000ffd70011fff00000ffcb000d0005ffe2fffa0045ffe90000000000eefff00006000e000000000025ffe90000ffdaffa8ffeaffc40000, 1024'hff8e000d0000000000310000ffedfff9000cfffffffcfff60001fffbffed006d00030009001cfffdfffc00000000ffd800000008fffcfff40015002500280008ffd3fffbffeffff3fff9ffda000400040000ffcb000ffffdffe1fffc0045fff30000000000f1fffb00000010000000000022fffb0000ffdbffa0fff5ffc60000, 1024'hff8f000c0000000000320000fff6fff3000c0001fffb000100010001fff2006b00020008001dfffdfffe00000000ffdc000000090002fffd0017002400270004ffda0000fff5fff4fff5ffdb000000000000ffcd000dfffdffdffffe0046fff40000000000ee0001ffff000c000000000023fff30000ffdcffa2fff3ffcb0000, 1024'hff8e000d0000000000320000fffdfff4000cfffffff9000400010002fff3006b00050005001dfffdfffe00000002ffe000000007000000020018002500280003ffe10002fffafff3fff9ffd70001fffc0000ffcb000d0000ffdefffe0045fff30000000000f1000100000007000000000023ffed0000ffdeffa5ffefffcc0000, 1024'hff8c000e0000000000320000fff7fff5000b0000ffffffff0001fff9ffec006d0006000c001bfffdfffb00000002ffdb00000007fffbfffe00190024002b0004ffdcfffefff6fff2fffcffd70003fffe0000ffc8000d0000ffdefffb0046fff20000000000f3fffd0002000e000000000024fff20000ffdeffa3ffeeffcb0000, 1024'hff8a000d0000000000340000fff7fff1000efffcfffcfffefffefff9fff0006e0005000e001cfffbfffb0000ffffffdc00000009fffdfffe001a0028002b0008ffd9fff8fff8fff2fff9ffdc0008fffc0000ffcb000dfffeffdcfffb0048fff50000000000f4fffa00050012000000000023fff20000ffd9ffa0fff1ffca0000, 1024'hff8b000c0000000000360000fff6fff3000efffffff7ffff0000ffffffee006f00080009001ffff9fffe00000002ffd9000000090000fffd00190026002c0004ffd9fffdfff7fff4fffaffd80006fffc0000ffcd000efffdffdcfffe0048fff20000000000f5fffd0002000c000000000022fff20000ffdcff9ffff2ffca0000, 1024'hff8c000c0000000000360000fff6fff6000f0001fff6fffc00000001ffed006f00070006001efff9ffff00000003ffda000000090003fffd00180026002c0004ffd9fffefff5fff4fff9ffd90005fffe0000ffcd0010fffeffdc00000048fff10000000000f4fffb0001000b000000000021fff20000ffdaff9ffff5ffcb0000, 1024'hff8c000c0000000000350000fff6fff7000d0001fff9fffdffff0000ffea006f00070006001dfffafffe00000005ffda000000090000fffe00190024002c0003ffdb0000fff5fff3fffbffd60003fffe0000ffcd00110001ffdd00010048ffee0000000000f4fffb0000000b000000000022fff10000ffdcffa0fff3ffcc0000, 1024'hff8b000c0000000000350000fff7fff5000efffdfffafffdfffdfffeffee006f00070008001cfffafffd00000003ffdb00000009fffefffe00190026002d0007ffdcfffcfff7fff4fffaffd90005fffd0000ffcd00110001ffdcffff0048fff00000000000f4fffb0002000e000000000022fff00000ffdbffa0fff3ffcc0000, 1024'hff8b000c0000000000360000fff6fff5000efffffff8fffdffff0000ffec006f00070007001efffafffe00000003ffda000000090000fffe00190026002d0005ffdafffefff6fff3fffaffd80005fffd0000ffcd0010ffffffdc00000048fff00000000000f5fffb0001000c000000000022fff10000ffdcff9ffff3ffcc0000, 1024'hff8c000e0000000000360000fff7fff2000dfffefff80001fffe0000fff1007000050006001cfff7fffd0000ffffffd8000000090001ffff0019002500300003ffdcfffefff7fff6fff8ffd80003fffc0000ffcb0010ffffffdbffff0048fff10000000000f6ffffffff000b000000000021fff00000ffdcffa1fff3ffd10000, 1024'hff89000f0000000000380000fffefff2000dffffffff0003fffdfff7ffe700720010000a001cfff9fffc0000fffeffd800000008fffd000e001d0021002e0003ffdffffcfffffff40000ffd7000bfff10000ffc80015fffcffdafffe0049fff10000000000f8fffb0002000d000000000028fff10000ffe5ffa2ffefffcd0000, 1024'hff85000d0000000000380000ffe7fff50010fffffff5ffeb0000fff0ffd8006e001b000d001dffe9fff90000ffffffca00000008fffdfff9001a00230034000dffc7ffe4ffef00060006ffd80017fff80000ffcb001d0003ffdb0001004dffea0000000000f2ffe30005001300000000001afffe0000ffdbff9a0000ffc70000, 1024'hff9100040000000000370000ffbe000b000dffffffe2ffc80009fff9ffb700650035000c002bffb6ffff00000021ff9f0000000c0003ffd500150022004b0019ffb4ffcdffca0032000bffd9001900160000ffe400230019ffd8000b004dffc40000000000cfffc50004001600000000ffff000f0000ffd8ff970018ffc40000, 1024'hffa0fffb00000000003c0000ffd700150017ffeaffc7ffb40004000fff96005c005500140040ffa1fffd0000003fffab00000014fffcfff10018002700530032ffcbffc1fff100270004ffdf003afff50000fffc0016002fffd5000d0052ffa60000000000a7ff99000a0015000000000002fff10000ffe7ffa60008ffc20000, 1024'hffa0fff700000000003e0000000b001a0025ffd5ffb0ffccfffd0008ffaa0068006500230042ffaefffe0000003effc000000013ffe8000c001b0029004000310009ffd10031ffff0021ffc20056ffba0000000100080023ffd7fff60055ffa900000000009dffa60012fffd000000000012ffbe0000fff4ffb1ffddffc10000, 1024'hff97fff900000000003c0000001200150026fffcffc9ffe1fff8ffe6ffc60074004a002c002effbbfffb0000002dffd700000011ffff0019001b002d002a00140004ffd30028fff00014ffca003cffc30000fff50003000bffd7ffe10053ffc00000000000afffcb001b001900000000001cffc50000ffd9ffa2ffd2ffbc0000, 1024'hff8bfffe00000000003d00000009ffff001c0001ffebfff8fff2ffeeffe300770020001d0020ffe2fffa00000015ffe20000001000060019001e002f0021000cfff1ffe3000fffedfffeffd9001cffe20000ffeb000f0008ffd4fff20054ffdb0000000000d4ffe80010001f000000000022ffda0000ffcdff94ffe3ffc00000, 1024'hff88000200000000003e0000fffefff30012fffcfff10005fffb0005fff20079000c00090023fff7fffd00000007ffdc0000000effff0009001d002a001f0007ffe8fffbfffefff00000ffd20008fff60000ffe400130008ffd2ffff0052ffea0000000000f1fffc00000009000000000022ffe00000ffd7ff8fffe8ffc10000, 1024'hffad000300000000003e0000ff850006001e0005ff8effb7003800a200070053ffdcff9b0066fff600360000fff2ffcc0000000d006effa0ffe5004c00190010ff7b0010ff950021ffd00008fff7005b00000006ffefffdeffe10036002700000000000000ccffe2ffc7ffc400000000fff1004f0000ffc0ff8c004fffbd0000, 1024'hff8f000700000000001d00000070ffb90025ffc50037003fff9eff700044004bfffc0064ffc5fff3ffcf0000ffdd003a0000000bffcc006a00420043001a00320032ff910061ffd8fff400170040ffa20000ffdb001b0010ffd5ffca004900240000000000a4ffed00670076000000000022ff9c0000ffa3ffc2ffd1ffee0000, 1024'hff8b000c00000000003a0000fffeffed0010fffefff80006fff50003fff1007200050001001bfffcffff0000fffeffdd0000000a0005000b001b0024002c0000ffde0000fffefff1fffaffdd0008fff50000ffd20017fffdffd900070048fff40000000000f7ffff0001000d000000000025ffef0000ffdbff9dfff6ffce0000, 1024'hff8e00020000000000390000ffcdffff0008000a0009ffe7fffeffe0ffd4006c0017000b0013fff1fffd00000006ffc000000008ffefffde001d00160030fffcffbefff0ffcf0005001bffcf000500120000ffdb002bfffcffd500060045ffeb0000000000dffff10008001700000000000f000d0000ffe3ff900008ffce0000, 1024'hff92fff000000000003e0000ffab000a0012000b0012ffb8ffe1ffbcffb7006a001700220004ffd0fff90000000fffa90000001afff8ffc80024000e00340011ffa3ffc3ffbd00130023ffec001d0016000000070050fffeffcd0012004effda00000000009fffc00018004700000000fffe001d0000ffc2ff820035ffd10000, 1024'hffa6ffe80000000000460000fff20002002bfff2ffd9ffceffba000effc300660026ffef0013ffbd000b00000020ffcc000000230022001d002000150029001affdbffcf0007000cfff6ffff0030ffde00000031005e0018ffce00410056ffbc000000000088ffb5000e002c00000000000affe80000ffc8ff870042ffd00000, 1024'hffaefff400000000004000000039fffc001fffddffc10013ffcd0048ffd6006b0044ffca0028ffd700150000002cffd9000000110005004f001d0008001e0003002b0014003c0000000fffc90024ffbc00000017004b002dffd500460050ffb80000000000baffe8fff7ffd8000000000023ffb000000007ffa10006ffc70000, 1024'hff96000800000000003500000027ffef0015ffe8ffdc0015ffe9001cffe900710029ffef0022ffec000300000010ffdf00000007fff4002c001b001900240006000e00080024fff70013ffcb001cffd30000ffdf0023001affdc0014004bffe00000000000f0fff20001ffee000000000029ffc00000fff1ffa6ffe7ffc00000, 1024'hff87000f0000000000320000fff2fffb000ffffeffeffff00002fffdffe00071001500050021ffeafffd00000007ffd000000006fffdfff8001600240031000affd5fff4fff4ffff0001ffd3000dfffb0000ffc500150005ffdfffff004affe80000000000feffed0003000a000000000020fff00000ffddff9efff7ffc00000, 1024'hff88000e0000000000330000ffe70002000e0000ffefffe50004fffcffd2006f001a000a0025ffdffffe00000011ffc5000000090003fff4001700250038000fffceffecffec0007fffcffd7001000010000ffcb00160008ffdf0002004cffdc0000000000f3ffe30002001000000000001dfffb0000ffdaff9fffffffc00000, 1024'hff8c000e00000000003400000000fffe0013fff7ffe6fff3fff90005ffd70072002200070024ffdfffff00000016ffcc0000000900010008001800240037000fffeafff2000400010004ffd6001affee0000ffd100160011ffde0004004cffd90000000000efffe300030009000000000022ffe40000ffdbffa6fff4ffc10000, 1024'hff8c001000000000003400000007fffe0013fffcffe7fff8fffa0004ffdf0074001b00020021ffe7fffe00000011ffd6000000070000000c0017002500320009ffecfff90007fff80002ffd20014ffed0000ffcb0014000dffdf0001004affe00000000000faffee00030006000000000025ffe10000ffdcffa5ffedffc00000, 1024'hff8900100000000000330000fff3fffe000d0001fff7fff50000fffbffe20074000e0006001dfff3fffc00000008ffd200000006fffdfffd0016002400300006ffdafffafff3fff8ffffffd30008fffe0000ffc600130005ffe0fffe0049ffe80000000000fefff50000000c000000000024fff50000ffdcff9ffff2ffc30000, 1024'hff8a000d0000000000340000ffe9fffa000b0000fffcfff30002fffbffe7007200060009001efff6fffb00000002ffd000000009fffffff500160025002c0009ffd0fff7ffeafffafffcffda000500070000ffcc00130002ffddfffe0049ffee0000000000f6fff5fffe0011000000000021fffd0000ffd8ff9cfff7ffc50000, 1024'hff8d000b0000000000360000fff6fff5000dfffefff9fffffffe0001ffeb007100090008001efff8fffd00000003ffd40000000a0000000100180023002a0006ffdcfffdfff6fff7fffcffd90006fffd0000ffd100130003ffdc0001004affee0000000000f1fffafffe000c000000000023fff20000ffdcff9efff3ffc90000, 1024'hff8c000b0000000000360000fffdfff3000efffdfff70003fffd0001fff0007100090006001dfff9fffd00000002ffdb00000009ffff00050019002400290004ffe0fffefffbfff5fffdffd70006fff90000ffcf00120003ffdb0000004afff10000000000f5fffc00010009000000000023ffec0000ffdcff9ffff0ffca0000, 1024'hff89000c0000000000360000fff7fff5000d0000fffc0000fffdfffbffec007300090009001bfffafffd00000003ffd700000009fffeffff001a0023002c0003ffddfffefff5fff50000ffd60005fffd0000ffcc00140001ffdbffff004afff00000000000f8fffc0001000d000000000023fff00000ffdaff9efff2ffcb0000, 1024'hff88000c0000000000370000fff7fff3000f0000fffcfffefff8fffbffed0073000600070019fff9fffd00000002ffda0000000a00010000001b0025002d0004ffdafffbfff5fff4fffcffdb0006fffd0000ffce00170001ffda0002004afff10000000000f9fff900030012000000000022fff00000ffd5ff9cfff7ffcb0000, 1024'hff89000c0000000000380000fff6fff4000ffffffffafffdfff80000ffeb007300070002001afffaffff00000003ffd80000000a0000ffff001b0023002e0003ffdafffffff5fff4fffcffd80005fffd0000ffcf001a0001ffda0007004affef0000000000fbfffb0001000d000000000022fff10000ffdaff9bfffaffcb0000, 1024'hff89000c0000000000380000fff5fff7000e0000fff9fff9fffc0000ffe9007200070002001cfff9fffd00000003ffd90000000affffffff001a0024002d0006ffd7fffdfff5fff4fff8ffd60004fffd0000ffce00190002ffdb0005004bffed0000000000fbfffaffff000c000000000022fff20000ffdcff9bfff8ffc90000, 1024'hff88000c0000000000370000fff4fff8000cfffefffcfffdfffefffdffea007400080007001cfff9fffc00000004ffd400000009fffcffff001a0024002d0006ffdcfffdfff4fff6fffcffd30003fffe0000ffce00160004ffdb0001004cffeb0000000000fafffcfffe000b000000000023fff20000ffddff9bfff3ffc90000, 1024'hff88000c0000000000380000fff5fff5000dfffffffbfffefffffffdffed007500070009001dfff7fffb00000002ffd50000000affff0000001a0027002c0007ffdcfffafff3fff7fffdffd7000400000000ffcf00130005ffd8fffe004cffee0000000000fafffbffff000e000000000022fff00000ffd8ff9afff0ffc90000, 1024'hff88000c00000000003a0000fff4fff4000d0000fffaffff00000000ffec007500070007001efffafffc00000001ffd50000000a00000000001a0026002d0005ffdafffdfff3fff6fffdffd60004ffff0000ffcf00130003ffd80000004cffef0000000000fbfffcfffd000b000000000022fff20000ffdaff9afff1ffcb0000, 1024'hff88000c00000000003a0000fff5fff6000c0002fffbffff0002ffffffec007400070009001dfffafffa00000006ffd70000000afffdfffd001b0029002f0006ffdcfffdfff0fff5fffaffd3000000040000ffce00110009ffd7fffe004dffec0000000000fdfffefffd000c00000000001fffee0000ffd7ff9affedffcc0000, 1024'hff84000d00000000003b0000fffbfff6000c0000000000010001fff8ffee00790003000d001c0000fff800000000ffdc0000000bfff80004001e0027002b0008ffe2fffffffaffecfffdffd00003fff90000ffcc00110002ffd7fff8004ffff00000000001010000fffd000b000000000027ffe90000ffdbff9bffe6ffca0000, 1024'hff7e000d00000000003b0000fff1fff500100006fffefffd0002fffaffec00780005000b001d0002fffc00000000ffdc000000090003ffff001c002e00290007ffdbfffafff0fff0ffffffd4000300010000ffcd00100001ffd7fffb004dffef000000000103fffdfffe0010000000000024fff10000ffd2ff93ffedffc70000, 1024'hff84000d00000000003a0000ffdbfff2000b0005fff6fff100070001ffe20071000a00050022ffe9fffd00000003ffc30000000a0005ffea0019002700390009ffc8fff1ffde000cffffffd70000000f0000ffd100160007ffd50004004bffe70000000000fbfff6fffb000e000000000017fffc0000ffd7ff93fffeffca0000, 1024'hff88000c00000000003d0000ffe7fff5000bfffcfff6fff1fffcfffbffd00070001d000a0025ffddfffd00000010ffbe0000000b00000000001f00220043000cffd6ffebfff0000c0006ffda0013fffb0000ffda001c0009ffd30008004affda0000000000ebffea0001001200000000001dfff90000ffe3ff9dfffbffcb0000, 1024'hff8b000a0000000000410000fff9fff50015fff6ffecffeffff4fff7ffcd00710026000e0022ffe0fff80000000cffc70000000bfff90011001f0027003c0013ffe0ffe40004fffc000bffda0026ffe60000ffdf001f000dffd30006004dffdb0000000000e5ffdd0006001500000000001effe90000ffe2ff99fff2ffc80000, 1024'hff8900060000000000410000fff6fff60012fffafff1fff4fff7fff3ffd20077001e00120022ffe7fff80000000cffc70000000dfff5000c002100240030000cffdcffeafffefff6000bffd3001fffec0000ffe2001e0009ffd300040053ffe00000000000edffe600070012000000000021ffed0000ffe0ff90ffefffbe0000, 1024'hff8400020000000000410000fff4fff30012fffafff7fffafff6fff4ffe4007d001000150021fff0fff700000006ffd000000010fff80007002000290025000dffdcffecfffbfff10004ffd60014fff30000ffe600190007ffd1fffd0056ffe70000000000f1ffef00050018000000000023ffea0000ffd5ff89ffebffbc0000, 1024'hff8300000000000000430000fff0fff00011fffdfff70001fffc0000fff2007e0006000d0024fff9fffc00000001ffd400000010ffff0001001e002b00200007ffd9fff7fff4fff1fffeffd50006fffd0000ffe700150001ffceffff0055ffee0000000000f7fffe00000010000000000022ffed0000ffd6ff84ffedffbf0000, 1024'hffac00000000000000440000ff82000000210004ff87ffb9003800ae000a0055ffdaff96006cfff7003a0000ffeeffca000000100077ffa2ffe5004f00170010ff750011ff930022ffcc000dfff9005c0000000efff0ffdaffdd003d002a00030000000000ceffe2ffc4ffc100000000fff000520000ffbeff840055ffbd0000, 1024'hff8b000700000000001f00000072ffb80025ffc100390042ff9dff6a004a004ffffa006affc3ffeeffcb0000ffdc00390000000cffca006d00440049001e00360033ff890061ffdbfff00017003fffa30000ffda00190015ffd2ffc5004e00230000000000abffed006a007b000000000020ff9a0000ff9dffbfffcdfff10000, 1024'hff89000b00000000003f0000fff3ffef000cfffffffa0005fffc0004fff1007700050003001ffffcfffd00000000ffd70000000b00020002001b002700320000ffd90000fff2fff5fffcffd9000300000000ffd300120000ffd40002004afff20000000000fd0002fffc000c000000000021fff50000ffdaff9afff0ffd20000, 1024'hff8c00080000000000400000ffdcfff9000d0007fffdfff00004fff2ffe00071000e0006001afff3fffd0000fff7ffc40000000bfffdfff1001a001e00340005ffc7fff5ffe10001000cffd3000600030000ffd50022fff7ffd500020049ffef0000000000eafff7fffb000d00000000001600010000ffe4ff94ffffffd90000, 1024'hff8d000100000000003e0000ffd30005000f000d0001ffdbfff5ffe6ffc6006f0016000a0013ffdffffd00000009ffb90000000f000cfff6001b001600350007ffbfffe1ffda00100010ffe0001100050000ffe700380004ffd50012004effdb0000000000cbffd90002001f000000000012000f0000ffd3ff920019ffd40000, 1024'hff98fffe00000000003c0000fff7fffc0014fff3ffecffebffdc000cffc8006f0025fff8001cffd8ffff0000001bffc5000000120009001b001b0018002e0012ffe3ffe5fffc000c0006ffe90022fff00000fffd003d0022ffd600260051ffcb0000000000c7ffceffff001700000000001bffef0000ffd6ff970012ffc30000, 1024'hff9a000300000000003b0000001affee0014ffe1ffde0010ffe2001effe400740028fff10024ffe600020000000fffce0000000dfff30029001c00160026000d00080002001ffffc0012ffd20021ffd50000fff2002d001bffd8001b004effda0000000000e1ffedfffbfff5000000000027ffc90000fff2ff9ffff0ffc00000, 1024'hff8b000c00000000003900000011ffec0013fffaffed0010fff30009fff300770011fffd001efff8000000000002ffdf0000000800000019001b00220025fffffff20004000efff00004ffd4000fffe70000ffd300180004ffd90006004bfff10000000000ff00010002000100000000002affdb0000ffe0ff9cffeaffc20000, 1024'hff8300100000000000370000fff4fff0000c0005fffc0002ffff0000ffec007500040001001dfffefffe0000fffeffd70000000700020000001a0025002b0000ffd40001fff0fff5fffbffd6000100010000ffc60016fffeffdc0004004afff400000000010c0001fffe000b000000000026fff50000ffdaff97fff5ffc30000, 1024'hff8200100000000000360000fff1fff3000b0000fffefffbfffffffeffe8007500040005001dfffbfffc00000001ffd200000008fffefffb001a0024002f0007ffd3fffdfff0fff8fffaffd7000300020000ffc600180002ffdc0004004cfff0000000000109fffbfffe000d000000000026fff60000ffdaff99fff8ffc20000, 1024'hff8300100000000000360000fffbfff6000efffffff7fffefffd0001ffe9007700080004001efff7fffd00000006ffd50000000800000003001a0027002e0007ffdffffefff8fff5fffbffd40006fffc0000ffc800160006ffdc0003004dffeb000000000109fffbffff000a000000000027ffec0000ffd8ff9afff2ffc10000, 1024'hff8300100000000000360000fff7fff5000c0000fffa0000ffff0002ffeb007800050003001ffffbfffd00000004ffd600000007ffff000100190027002d0004ffdc0001fff4fff4fffcffd4000200000000ffc700120004ffdc0001004bffee00000000010cfffefffe000a000000000028fff00000ffdaff99ffefffc10000, 1024'hff83000f0000000000370000ffeefff3000c0000fffdfffb0002fffdffeb007600040008001efffcfffc0000ffffffd200000008fffdfff700190027002f0006ffd3fffdffedfff6fffdffd6000200050000ffc600120000ffdaffff004bfff2000000000108fffdffff000e000000000024fff60000ffdaff97fff3ffc60000, 1024'hff85000c0000000000390000ffecfff4000d0000fffafff80001fffdffe80074000600090020fff6fffd00000001ffd10000000a0001fff8001a002700300006ffcefff9ffedfff8fffaffd9000500030000ffcc0013fffeffd90001004cfff00000000000fffff700010010000000000021fff90000ffd9ff97fff8ffc80000, 1024'hff87000b00000000003a0000fff4fff5000efffefff7fffbfffdffffffe70075000b00080020fff6fffd00000005ffd40000000bffffffff001b0025002f0006ffd8fffbfff6fff5fffcffd60009fffb0000ffd000150001ffd90002004dffec0000000000fbfff80000000d000000000023fff20000ffdbff9afff4ffc80000, 1024'hff87000b00000000003a0000fff7fff4000ffffefff7fffffffcffffffeb0075000b0007001ffff7fffd00000003ffd70000000affff0003001b0027002d0006ffdcfffbfff8fff4fffcffd60008fff90000ffd100140001ffd90000004cffed0000000000fbfffa0000000d000000000023ffee0000ffdbff99fff1ffc80000, 1024'hff86000c00000000003a0000fff6fff5000e0001fffafffefffffffdffeb007600070008001dfff9fffc00000002ffd50000000affff0000001b0026002d0005ffdbfffdfff5fff4fffdffd40004fffd0000ffce00150002ffd80000004dffee0000000000fefffdffff000c000000000023ffef0000ffdaff98fff1ffc90000, 1024'hff85000c00000000003a0000fff6fff6000e0002fffbfffefffefffdffeb007700060007001cfff9fffc00000003ffd60000000a00010002001b0027002d0005ffdbfffcfff3fff5fffcffd50003ffff0000ffce00160004ffd80001004effed000000000100fffcffff000d000000000023fff00000ffd7ff97fff2ffc90000, 1024'hff85000c00000000003a0000fff4fff7000d0001fffbfffdffff0000ffea007800060005001dfffafffc00000003ffd40000000a00000000001a0026002d0006ffdbfffefff1fff6fffeffd4000200010000ffce00170006ffd80002004effec000000000101fffbfffc000b000000000023fff00000ffd8ff97fff2ffc90000, 1024'hff84000b00000000003a0000fff2fff6000b0000fffffffdfffffffdffe9007800050008001efffdfffa00000003ffd60000000afffc0000001b0026002b0006ffd8fffdfff1fff3fffdffd4000200010000ffcf00150005ffd80000004effed000000000101fffbfffd000e000000000025fff30000ffdaff96ffefffc60000, 1024'hff83000a00000000003b0000fff1fff2000dfffdfffefffffffffffbffee00780005000d001efffdfffa00000000ffd40000000bfffafffc001c0029002b0009ffd9fffafff1fff3fffeffd5000400010000ffd100130003ffd6fffd004ffff0000000000100fffdffff0010000000000023fff00000ffd8ff93ffeeffc70000, 1024'hff83000900000000003d0000fff2fff1000e0001fffb00000000fffeffef00780003000b0020fffbfffc00000001ffd70000000c0000fffd001d002a002b0005ffd7fffcfff1fff2fffbffd6000200010000ffd300110000ffd4fffe004ffff1000000000100fffe0000000f000000000022ffef0000ffd6ff92ffefffc80000, 1024'hff83000900000000003e0000fff2fff3000f0001fffafffe00000000ffed0078000400090020fffdfffd00000002ffd80000000c0000fffd001d002a002c0005ffd8fffefff2fff0fffbffd4000200000000ffd300120000ffd40000004fffef000000000100fffeffff000d000000000022ffef0000ffd8ff92fff0ffca0000, 1024'hff82000800000000003e0000fff2fff6000e0003fffdfffc0001fffbffea00780005000c001ffffefffb00000005ffd90000000cfffcfffc001e002a002b0006ffd8fffdfff1ffeefffcffd1000100010000ffd300130002ffd4fffe0050ffed000000000100fffe0000000f000000000022ffee0000ffd8ff91ffedffc80000, 1024'hff7f000600000000003e0000fff2fff4000e00000003fffffffcfff7fff0007cfffc0010001d0006fffa00000002ffdd0000000dfffafffd001f002b00250006ffd9fffefff3ffe6fffcffd4000100000000ffd70012fffeffd4fffc0051fff2000000000101000000020014000000000027ffef0000ffd4ff8dffebffc40000, 1024'hff81000500000000003f0000ffeffff000100002ffff0000fffffffefffa007cfff6000a001e0007fffc0000fff7ffde0000000e0001fffb001c002c001f0004ffd40000fff0ffe7fff6ffd6fffb00030000ffd80012fff8ffd2fffd0051fff80000000001010007fffe0011000000000025fff00000ffd5ff87ffefffc70000, 1024'hff8300060000000000400000ffe9ffed000900060002000900060003fffb0078fff8000700200003fffd0000fffbffd70000000d0003fff7001e002b0026fffdffd10004ffe4fff3fff3ffd2fff0000f0000ffd70010fffdffcf00000050fff50000000001020010fff9000b00000000001efff60000ffd8ff8afff0ffcf0000, 1024'hff8500080000000000430000ffedffea0008ffff0007000d0002fffcfffd007bfff8000d001c0002fff90000fff8ffd30000000efffbfffa00210029002e0000ffd90002ffeafff3fffcffd4fff600090000ffd80010ffffffcbfffb004ffff80000000000fe000efffa000d00000000001efff20000ffd9ff91ffeaffd70000, 1024'hff8200080000000000480000fff0ffe8000e000400070008fffffff6fff3007affff0011001b0007fff80000fff7ffdc0000000ffffd00040024002d002f0002ffd6fffbfff0ffebfffdffd7000000000000ffd80010fffcffcafffb0050fff80000000000fe0007ffff0015000000000020fff30000ffd8ff8effe8ffd90000, 1024'hff7d00050000000000490000ffebffe8000e000000080003fffdfff2ffef007c00000014001c000afff70000fff6ffd80000000ffff8ffff0024002a002c0005ffcffff8fff1ffea0001ffd60006fffc0000ffdb0016fff9ffcbfffd0053fff90000000000fe000100000016000000000022fff70000ffd9ff89ffedffd10000, 1024'hff7d00010000000000480000ffe7ffea000e000100060000fffafff1ffef007ffffe0015001e0003fff70000fffaffd500000011fffafffd0024002b00250004ffccfff4ffedffeafffdffd7000500000000ffe40018fffaffcafffe0056fff50000000000fc00000002001b000000000022fff80000ffd4ff80ffefffc60000, 1024'hff80fffe00000000004a0000ffe9ffe60013fffcfffc0005fffa0000fff5007f0001000f0023fffefffe0000fff8ffd0000000130001ffff0023002d00230006ffd1fff7ffeefff0fffeffda000500000000ffec0018fffaffc700040057fff50000000000f900000001001400000000001ffff10000ffd6ff7bfff4ffc80000, 1024'hffabfffe00000000004b0000ff84fffa00250003ff7effb9003500ba000b0056ffd9ff8e0070fff8003e0000ffedffce00000013007fffa4ffe700500019000dff700014ff970020ffc90010fffd005800000014fff3ffd7ffd80047002c00060000000000d1ffe0ffc4ffbc00000000ffee00520000ffbcff81005dffc00000, 1024'hffaf000700000000001000000056ff850036000e005a0048ff39ff9a00560026ffa1fffdff85005800000000ffd2008b0000000dfffd002e00490017fffaffd9001afff70033ff88fffb00590013ffd1000000060063ffd4ffdf0032fffd00670000000000850021006b009d00000000001eff9d0000ff74ffb8003cfff50000, 1024'hffaf00090000000000210000fffdffac001f0016004e001dff69000200310026ff83ff94ffab007a00360000ffe2004a0000000d0000ffd50048fff4000dffb1ffd10064ffe9ff8cffd20012ffc0001b000000010094ffaaffde009cfffc00480000000000d4006e0035003300000000001bfff70000ffdeff8f009bfff10000, 1024'hffaf00080000000000220000fff7ffad00200017004d0014ff6cffff00290024ff87ff97ffad007900350000ffde00490000000f0001ffd50047fff1000dffb6ffc9005dffeaff8fffd30013ffc60016000000010095ffa6ffe0009bfffe00470000000000cd00670034003400000000001cfffe0000ffe2ff90009efff30000, 1024'hffae00060000000000200000fff7ffb0001f0014004b0013ff6afffd00220023ff94ff99ffb0007100350000ffe300430000000d0003ffdb0045ffee000cffb8ffcc0056ffeeff98ffd80014ffce000f000000050099ffa9ffe2009bfffe003f0000000000c1005e0033003500000000001d00000000ffe4ff9300a0ffee0000, 1024'hffb2000600000000001e00000002ffad001f000f0047001bff63000100230025ff96ff99ffb1006b00340000ffe9003f0000000d0002ffe50045ffee0008ffb8ffd70056fff5ff98ffdb0018ffd4000c0000000c009affb2ffe2009efffe003d0000000000c0005c00350036000000000020fff80000ffe0ff93009bffe30000, 1024'hffb4000800000000001e00000010ffa40020000d0046002aff5f000600310028ff8fff95ffae007400340000ffe200480000000dfffeffed0046ffed0003ffb3ffe20060ffffff8fffda0016ffd10006000000090097ffb0ffe2009dfffe00470000000000cc006a00350030000000000025ffec0000ffe2ff930092ffe30000, 1024'hffaf000a00000000001e0000000bffa3001d0013004e002eff670005003c0028ff82ff93ffad008100340000ffd900500000000b0000ffe70045fff10000ffafffd90067fff7ff8affd20014ffc3000f0000ffff0091ffa7ffe30098fffc00510000000000d900770032002f000000000026fff30000ffe2ff910090ffe70000, 1024'hffab000c00000000001d00000000ffa3001900170057002bff6e0001003c0028ff7aff96ffac008900330000ffd4004d0000000a0000ffdd0044fff00001ffaeffce0069ffecff8bffd00014ffbc00190000fff7008fffa2ffe40096fffc00560000000000df007b002f0030000000000027ffff0000ffe2ff900093ffe90000, 1024'hffa9000c00000000001c00000000ffa200180017005a002cff6dfffe003b0028ff7aff99ffac008900320000ffd5004d0000000a0000ffde0045fff10000ffafffce0067ffebff8bffd10016ffbd001a0000fff7008fffa3ffe40095fffc00560000000000df007900300034000000000028ffff0000ffdfff900092ffe70000, 1024'hffa9000c00000000001c00000002ffa0001900150058002dff6b0000003d0028ff79ff98ffac008900320000ffd5004e0000000affffffde0045fff20000ffb0ffcf0067ffedff8affd00017ffbe00190000fff8008fffa4ffe40096fffc00570000000000e1007900310034000000000028fffc0000ffdeff8f0092ffe50000, 1024'hffaa000c00000000001c0000ffffffa1001900160057002bff6d0000003d0028ff79ff97ffac008700330000ffd4004c0000000affffffda0045fff10001ffaeffcd0068ffeaff8bffd00015ffbc001b0000fff7008fffa2ffe30096fffc00570000000000e1007a00310032000000000026fffd0000ffe0ff8e0094ffe70000, 1024'hffaa000c00000000001d0000fffcffa30019001800570028ff6efffe003a0027ff7bff98ffac008300330000ffd6004a0000000b0001ffd80046fff20004ffafffcb0065ffe7ff8effd00015ffbc001d0000fff80090ffa3ffe20096fffc00540000000000de007800310034000000000023ffff0000ffdeff8f0096ffea0000, 1024'hffab000c00000000001e0000fffcffa4001a001700550025ff6cffff00350026ff80ff97ffac008000330000ffd900490000000b0001ffda0046fff10008ffb1ffcc0062ffe9ff91ffd10016ffc0001a0000fffa0092ffa6ffe20098fffc00500000000000da007300310034000000000022ffff0000ffdfff910098ffeb0000, 1024'hffac000b00000000001e0000ffffffa7001b001500540024ff6affff00320027ff82ff98ffac008000330000ffdd00480000000bffffffdc0046fff10007ffb2ffd10063ffecff8effd50015ffc300180000fffd0093ffa9ffe20099fffc004d0000000000d7007000320034000000000023fffc0000ffdfff910096ffe90000, 1024'hffad000a00000000001e00000001ffa5001d001500520024ff68ffff00340027ff81ff98ffab008000330000ffdb004b0000000cffffffdd0046fff10005ffb2ffd10062ffeeff8cffd40016ffc400160000fffe0093ffa8ffe20099fffd004f0000000000d7007000340035000000000023fff90000ffdeff8f0096ffe90000, 1024'hffab000900000000001e00000001ffa5001c001500540026ff68ffff00350027ff81ff98ffac008200340000ffdc004d0000000cffffffdd0047fff10004ffb1ffd10064ffeeff8bffd30015ffc200160000fffe0093ffa6ffe20099fffd004f0000000000d8007200340035000000000024fff90000ffdfff8f0096ffe90000, 1024'hffaa000900000000001e00000001ffa4001d001400530025ff67ffff00360027ff80ff98ffac008200340000ffdb004e0000000cffffffdc0047fff20004ffb2ffd00063ffefff8affd20016ffc300150000fffe0093ffa5ffe20099fffd00500000000000d9007100350036000000000024fff80000ffdeff8e0097ffe80000, 1024'hffaa000900000000001e00000000ffa5001d001500520024ff68000000350027ff80ff97ffad008100350000ffdc004d0000000c0000ffdb0047fff20004ffb1ffcf0064ffeeff8affd10015ffc200160000fffe0093ffa4ffe2009afffd004f0000000000da007200350035000000000024fff90000ffdfff8d0098ffe70000, 1024'hffaa000800000000001e0000ffffffa5001d001500550024ff66fffc00340028ff81ff99ffab008200350000ffdc004c0000000cfffeffda0048fff00003ffafffcf0064ffedff89ffd50015ffc300160000ffff0095ffa3ffe1009afffd00500000000000d8007100370037000000000024fffa0000ffdfff8c0099ffe70000, 1024'hffaa000700000000001f0000ffffffa3001f001500540023ff62fffb00360028ff7fff99ffa9008000350000ffdb004d0000000e0000ffd90049fff10003ffb0ffcd0061ffedff89ffd30018ffc40016000000020098ffa3ffe0009cfffe00510000000000d700700039003b000000000022fff90000ffdaff8a009dffe80000, 1024'hffab000600000000002000000000ffa4001f001500530024ff60ffff00360028ff80ff94ffa9008000370000ffdd004e0000000e0001ffdb0049ffef0004ffaeffce0064ffeeff8affd10017ffc2001500000004009bffa3ffe000a0fffe004f0000000000d7007200380038000000000022fff90000ffddff8a00a0ffe90000, 1024'hffab000600000000002000000000ffa5001f001400530023ff60000000350028ff80ff93ffa9008100370000ffdd004e0000000e0000ffdb0049ffef0004ffafffcf0065ffeeff89ffd20016ffc2001500000004009cffa4ffe000a1fffe004e0000000000d7007100370037000000000022fff80000ffdeff8a00a0ffea0000, 1024'hffaa000500000000002000000000ffa5001f001400560023ff5efffc00330029ff81ff95ffa8008300370000ffdd004e0000000efffeffdc004affed0002ffaeffcf0065ffefff87ffd60016ffc4001300000005009effa2ffe000a1fffe004f0000000000d6007000390039000000000024fff90000ffdfff8900a0ffe80000, 1024'hffaa00030000000000200000fffeffa30021001300570021ff59fff90035002aff7fff96ffa5008300370000ffda004e0000000fffffffda004affecffffffadffcb0062ffeeff86ffd6001affc600130000000800a2ffa0ffdf00a3ffff00520000000000d3006d003c003e000000000023fffb0000ffdbff8500a6ffe70000, 1024'hffac00010000000000210000fffdffa10021001200530022ff58000000360028ff80ff92ffa8007f00390000ffdd004e000000110001ffd9004bffedffffffadffc80062ffecff89ffd0001bffc400160000000d00a3ffa2ffde00a8000000500000000000d3006e003c003d000000000020fffb0000ffdbff8300aaffe60000, 1024'hffad00000000000000220000ffffffa30021001000500024ff59000200370027ff84ff92ffa8007d003a0000ffe3004d00000011fffcffd4004cffed0005ffaeffcf0065ffedff8bffd30015ffc200160000000e00a2ffa6ffdd00a70000004c0000000000d20071003c003800000000001cfff30000ffddff8600a7ffeb0000, 1024'hffac000000000000002300000000ffa8002400140050001eff58fffd00340027ff83ff95ffa5007a003a0000ffe8005200000012fffeffd2004efff1000bffafffd20063ffecff87ffd20015ffc100170000000d00a0ffa7ffdb00a4000000480000000000d0006d0040003d000000000019ffed0000ffd7ff8700a6fff20000, 1024'hffaa000000000000002500000003ffab002700140053001aff53fffa0031002aff81ff94ffa20080003b0000ffe6005800000013ffffffd70050fff0000affaeffd50066fff2ff7dffd40015ffc400100000000d00a4ffa2ffda00a6000000480000000000cf006a0041003f00000000001dffec0000ffd8ff8700a8fff60000, 1024'hffa8ffff00000000002600000002ffa8002900150056001aff4dfff70030002bff82ff92ff9f0085003c0000ffe2005a000000130000ffda0051ffee0005ffabffd10065fff3ff7affd60017ffc7000d0000000f00abff9effda00ab0000004b0000000000d0006a0043004300000000001ffff10000ffd8ff8200aefff30000, 1024'hffa8fffc0000000000260000fffcffa3002800130059001bff47fff60031002bff81ff91ff9d0084003d0000ffe2005400000014fffeffd40052ffea0003ffa9ffc90063ffedff7fffd7001bffc700120000001500b3ff9effd900b20001004e0000000000d0006a0046004700000000001dfff70000ffd6ff7c00b8ffed0000, 1024'hffaafffc0000000000270000ffffff9e002a000f004f001bff4300000035002aff80ff89ffa0007b003f0000ffdf0054000000170003ffd70052ffe90005ffacffc80061fff3ff84ffce001effc9000c0000001900b7ff9dffd900b80003004d0000000000d1006a0044004300000000001cfff20000ffd7ff7c00bfffed0000, 1024'hffd6fffd0000000000270000ffaeffd20027ffffffe6ffb8ffaf008000320000ff74ff44fff2003800420000ffc20039000000130041ffad00130012000cffe4ff580040ffc4ffc9ff570027ffab003c00000018007bffa6ffed00ba0000002c0000000000a700340001fffb00000000ffed004100000005ff8000e5fff30000 };

wire [47:0] airplane4_image [1023:0] = { 48'h1100120014, 48'h1100130014, 48'h1200130015, 48'h1200130015, 48'h1300140015, 48'h1200130015, 48'h1200130015, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1400150016, 48'h1400150016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1200130015, 48'h1200130015, 48'h1100120014, 48'h1100120014, 48'h1100120014, 48'h1100110014, 48'h1000110014, 48'h1000100013, 48'hf000f0012, 48'he000f0011, 48'he000e0011, 48'hd000e0011, 48'he000f0011, 48'h1100120014, 48'h1100130014, 48'h1200130015, 48'h1300130015, 48'h1300140015, 48'hf00100011, 48'hd000e000f, 48'h1200130015, 48'h1400150016, 48'h1300140015, 48'h1300140016, 48'h1300140015, 48'h1300140015, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140016, 48'h1300140015, 48'h1200130015, 48'h1200130015, 48'h1100120014, 48'h1100120014, 48'h1100110014, 48'h1000110014, 48'h1000100013, 48'hf00100013, 48'hf00100013, 48'he000f0012, 48'he000f0011, 48'hd000e0011, 48'he000f0011, 48'h1100120014, 48'h1100130014, 48'h1100130014, 48'h1300140016, 48'h9000b000f, 48'h600090009, 48'h500050008, 48'h600060009, 48'h1000120013, 48'h1400150016, 48'h1300140015, 48'h1300140015, 48'h1200140015, 48'h1300150015, 48'h1300140015, 48'h1300140015, 48'h1300140015, 48'h1300140015, 48'h1200130015, 48'h1200130015, 48'h1100130015, 48'h1100120014, 48'h1100120014, 48'h1100110014, 48'h1000110014, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'he000e0012, 48'hd000e0011, 48'hd000e0010, 48'he000f0012, 48'h1100120014, 48'h1100130014, 48'h1100120014, 48'h1200140015, 48'hfffe00020008, 48'hfff7fff90001, 48'h400040008, 48'h100020004, 48'h200040004, 48'hf000f0010, 48'h1400140015, 48'h1200140015, 48'h1100140014, 48'h1200150015, 48'h1000120013, 48'hf00100011, 48'h1200130015, 48'h1200130015, 48'h1100130014, 48'h1100120015, 48'h1100120015, 48'h1100120015, 48'h1100110014, 48'h1000110014, 48'h1000100013, 48'h1000100013, 48'hf00100013, 48'hf00100013, 48'he000e0013, 48'he000e0011, 48'hd000f0010, 48'he000f0011, 48'h1100120014, 48'h1100130014, 48'h1100120014, 48'h1100130014, 48'hc000d0013, 48'hfff5fff60005, 48'hfff4fff80000, 48'h60004, 48'hffff00020001, 48'hffff00000000, 48'hc000d000d, 48'h1300150015, 48'h1100130015, 48'h1200140016, 48'h1100120014, 48'h9000a000b, 48'h1300140016, 48'h1300140015, 48'h1200130015, 48'h1100120015, 48'h1100120015, 48'h1100110014, 48'h1000110014, 48'h1000100013, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'he000f0012, 48'he000f0010, 48'hd000f000f, 48'he000f0011, 48'h1100120014, 48'h1100120014, 48'h1100120014, 48'h1100120014, 48'h1300130016, 48'h8000c0012, 48'hffedfff30000, 48'hfff4fffa0000, 48'h100030007, 48'h3, 48'hfffcfffdfffd, 48'h8000a000a, 48'h1400150017, 48'h1100110015, 48'h200030005, 48'hfff5fff7fff9, 48'h300040006, 48'h1000110013, 48'h1100120014, 48'h1100110014, 48'h1100120015, 48'h1100110014, 48'h1000110014, 48'h1000110014, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'he000f0011, 48'hd000e0010, 48'hd000e0010, 48'he000f0010, 48'h1000110013, 48'h1100120014, 48'h1100120014, 48'h1100120014, 48'h1200120013, 48'h1000140013, 48'h4000a000f, 48'hfff0fff20003, 48'hfff6fff70003, 48'h20006, 48'hfffe00000001, 48'hfffbfffdfffd, 48'h200030004, 48'hfffbfffbffff, 48'hfff3fff3fff7, 48'hffebffebffee, 48'hfff9fff9fffc, 48'h1000100014, 48'hd000e0010, 48'he000f0012, 48'h1200130015, 48'h1100110014, 48'h1000110014, 48'h1000110014, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'he000f0012, 48'hd000e0010, 48'hd000e0011, 48'he000e0012, 48'hd000e0011, 48'h1000110013, 48'h1000110013, 48'h1000110013, 48'h1100120014, 48'h1200130014, 48'h1200120014, 48'h1100130014, 48'h400060010, 48'hffeefff10000, 48'hfff7fff80002, 48'hfffe00000003, 48'hfffe0000ffff, 48'hfff5fff6fff6, 48'hffedffedffef, 48'hfffafffafffd, 48'hfffafffbfffe, 48'hffffffff0003, 48'h1400140017, 48'hd000d0010, 48'ha000a000d, 48'h1000110013, 48'h1000110014, 48'h1000110014, 48'h1000110014, 48'h1000100013, 48'hf00100013, 48'hf00100013, 48'hf00100013, 48'he000e0011, 48'hb000b0011, 48'h900090010, 48'hc000c0011, 48'hf00110013, 48'h1000110013, 48'h1000110013, 48'h1000110013, 48'h1100110014, 48'h1300110015, 48'h1300110014, 48'h1100150015, 48'h3000c, 48'hfff1fff1fffb, 48'hfffeffff0003, 48'hfffcfffefffd, 48'hfff7fff8fff7, 48'hfff9fff9fffa, 48'hfffbfffcffff, 48'h70008000a, 48'h100020005, 48'hc000c000f, 48'hfff6fff6fffa, 48'hfff2fff2fff7, 48'h60007000a, 48'h1100130014, 48'h1000110013, 48'h1000110013, 48'hf00100013, 48'h1000100013, 48'hf00100013, 48'ha000a000e, 48'hfffefffe0003, 48'hffefffeffff7, 48'hffe7ffe7fff1, 48'h100010009, 48'hf00100011, 48'hf00110011, 48'hf00110012, 48'h1000120013, 48'h1000120013, 48'h1100120013, 48'h1100120013, 48'h1100120013, 48'h1100120014, 48'h300040007, 48'hfffcfffdffff, 48'hfffbfffdfffd, 48'hfffafffcfffb, 48'hfffeffffffff, 48'hfffafffbfffd, 48'hfffcfffdffff, 48'h100020004, 48'hfffafffbfffd, 48'hffeeffeefff3, 48'hffedffedfff2, 48'ha000b000d, 48'h1100120012, 48'h1000110012, 48'h1000110012, 48'hf00100012, 48'hb000c000f, 48'h10005, 48'hfff0fff1fff5, 48'hffe5ffe6ffe9, 48'hffd9ffdbffe1, 48'hffdeffe0ffe9, 48'h30005000b, 48'he000f000f, 48'he000f0010, 48'hf00100010, 48'hf00110011, 48'h1000110011, 48'h1000110011, 48'h1100110012, 48'h1100120012, 48'h1100110012, 48'hf00100011, 48'h10002, 48'hfff8fff9fffa, 48'hfffdfffffffe, 48'hfffeffffffff, 48'hffff00000002, 48'hfffcfffdffff, 48'hfff4fff5fff7, 48'hfff5fff6fff8, 48'h100010004, 48'hfff9fff9fffd, 48'h9000a000b, 48'h1000110012, 48'hf00100013, 48'he000f0011, 48'h200040006, 48'hfff3fff5fff8, 48'hffe9ffebffed, 48'hffe3ffe4ffe7, 48'hffdaffdcffdb, 48'hffd1ffd3ffd4, 48'hffeffff2fff5, 48'hc000e000f, 48'he000e000e, 48'he000e000e, 48'hf000f000f, 48'hf000f000f, 48'hf000f000f, 48'h1000100010, 48'h1100110011, 48'h1100110011, 48'h1000100011, 48'h1000110011, 48'hf00100010, 48'hffff00010000, 48'hfff9fffafffa, 48'hfffeffffffff, 48'h400050006, 48'hffff00000002, 48'hfffcfffdfffe, 48'hfff7fff7fff9, 48'h100020003, 48'h600070008, 48'h80009000b, 48'hf00100013, 48'h90009000e, 48'hfff7fff9fffc, 48'hffe5ffe9ffea, 48'hffe7ffeaffeb, 48'hfff1fff4fff5, 48'hfffcfffeffff, 48'hffeeffefffee, 48'hffedffeeffee, 48'h700070009, 48'ha000b000b, 48'he000d000d, 48'he000d000d, 48'hf000e000e, 48'hf000e000e, 48'hf000e000e, 48'hf000f000e, 48'h10000f000f, 48'h10000f000f, 48'h100010000f, 48'hf0010000f, 48'h100010000f, 48'hb000c000c, 48'hfffdfffefffd, 48'hfffafffbfffc, 48'hffff00000002, 48'hfffcfffdfffe, 48'hfffeffff0001, 48'hfffeffff0000, 48'hfff8fff9fff9, 48'h700080009, 48'ha000a000d, 48'h4, 48'hfff1fff2fff5, 48'hffe9ffecffee, 48'hfff3fff6fff8, 48'h300050006, 48'h9000a000b, 48'h400040004, 48'hfffcfffbfffc, 48'h800050007, 48'hb0008000a, 48'ha0008000a, 48'hd000b000a, 48'hd000b000b, 48'he000c000b, 48'he000c000c, 48'he000d000c, 48'he000d000d, 48'hf000e000d, 48'hf000e000d, 48'he000e000d, 48'he000f000c, 48'he000e000c, 48'he000e000e, 48'h900090009, 48'hfffafffafffc, 48'hfff9fff9fffb, 48'hfffeffff0000, 48'h100020004, 48'h300040006, 48'hfff8fff9fffa, 48'hfff7fff8fff9, 48'hfff2fff2fff6, 48'hffebffebffef, 48'hfff3fff4fff7, 48'h300040006, 48'hb000d000f, 48'h80009000a, 48'hffffffff, 48'hfffefffe, 48'h700050006, 48'hb00070008, 48'hb00060006, 48'hb00070007, 48'hb00090008, 48'hb000a0008, 48'hc000a0009, 48'hc000a000a, 48'hd000b000a, 48'hd000c000a, 48'hd000d000b, 48'hd000d000b, 48'hd000d000b, 48'hd000d000a, 48'hd000d000a, 48'hc000c000a, 48'hd000c000b, 48'h600060006, 48'hfffcfffdffff, 48'h200030004, 48'h100020004, 48'hfff5fff5fff7, 48'hffe9ffebffec, 48'hffe8ffe9ffeb, 48'hffe9ffe9ffed, 48'hfffafffafffe, 48'he00100011, 48'hd000e000e, 48'hffffffff0001, 48'hfffafff9fffa, 48'h500030000, 48'hb00080006, 48'ha00070005, 48'h900060003, 48'ha00050002, 48'ha00060004, 48'ha00080004, 48'hb00090005, 48'hb00090006, 48'hb00090007, 48'hd00090006, 48'hc000a0006, 48'hb000b0008, 48'hc000b0008, 48'hd000b0008, 48'he000a0008, 48'hd000a0008, 48'hc000a0008, 48'hb00090008, 48'h900080008, 48'hfff9fff9fffc, 48'hfff2fff3fff5, 48'hffe9ffebffed, 48'hffe6ffe7ffe9, 48'hffe9ffebffec, 48'hfff9fffafffc, 48'h80007000b, 48'hc000c000f, 48'h200050006, 48'hfffcfffffffd, 48'hfffdfffcffff, 48'hfffbfffcfffe, 48'h40004ffff, 48'h900050002, 48'h800040001, 48'h800040000, 48'h700040000, 48'h800050001, 48'ha00060000, 48'hb00070001, 48'hb00070002, 48'hc00070003, 48'hc00070003, 48'hb00080004, 48'hb00090004, 48'hd00090004, 48'he00090004, 48'he00090004, 48'hc00080004, 48'ha00080005, 48'h900080008, 48'h600060007, 48'hffeffff0fff3, 48'hffdfffe0ffe3, 48'hffe3ffe5ffe8, 48'hfff2fff4fff8, 48'h300060009, 48'hc000e0010, 48'h80007000b, 48'hfffcfffbfffd, 48'hfff6fff8fff7, 48'h100040004, 48'hfff9fffbffff, 48'hffeaffebffed, 48'hfffcfffcfff8, 48'h800040000, 48'h70002fffe, 48'h70003fffd, 48'h60002fffc, 48'h70002fffd, 48'hb0004fffd, 48'ha0005ffff, 48'hb0005ffff, 48'hd0005fffe, 48'hb00050000, 48'hb00050000, 48'hb0006ffff, 48'he00070000, 48'he00060000, 48'hc00060000, 48'hb00070003, 48'h900060005, 48'h1, 48'hfff3fff4fff7, 48'hffe6ffe8ffeb, 48'hffe9ffebffee, 48'hfffe00010004, 48'he00100014, 48'ha000d000f, 48'hfffcfffd0000, 48'hfffafffafffd, 48'hfffefffeffff, 48'hfff8fff9fff7, 48'hfff9fffafffa, 48'hfff8fff8fff9, 48'hfff1ffefffed, 48'hfff9fff6fff1, 48'h70002fffa, 48'h60001fff9, 48'h60001fff9, 48'h60000fff8, 48'h60001fff9, 48'h80001fffb, 48'h70002fffe, 48'h80003fffd, 48'hb0004fffc, 48'hb0004fffd, 48'hb0004fffc, 48'hc0005fffb, 48'hb0005fffd, 48'hb0004ffff, 48'h900050001, 48'h40001fffe, 48'hfff8fff7fff7, 48'hffedffedffef, 48'hffeefff0fff2, 48'hfffbfffdfffe, 48'h9000a000b, 48'hd000d000d, 48'h500040002, 48'hfffafff9fff8, 48'hfffdfffcfffd, 48'h500060008, 48'h600070008, 48'hfffbfffcfffb, 48'hfff9fff8fff6, 48'hfffdfffbfff6, 48'h2fffdfff7, 48'hfff9fff3ffee, 48'h2fffcfff3, 48'h70000fff6, 48'h6fffffff4, 48'h6fffffff4, 48'h70000fff5, 48'h1fffcfff9, 48'h400000000, 48'h40001fffe, 48'h70001fffa, 48'ha0002fff9, 48'hb0003fff8, 48'hb0003fff7, 48'h90003fffb, 48'h40001fffd, 48'hfff8fff7fff7, 48'hffeeffedffee, 48'hffedffeeffef, 48'hfff5fff6fff9, 48'h500070009, 48'hb000d000e, 48'h500050003, 48'h2fffefff9, 48'h3fffefff5, 48'h1fffcfff5, 48'hfffefffbfff9, 48'h10001, 48'hfffe00000001, 48'hfffeffff0000, 48'hfffcfffafffb, 48'hfffcfffafff4, 48'h40000fffa, 48'hfffcfff8fff7, 48'hfff6fff3ffef, 48'h4fffdfff1, 48'h6fffefff1, 48'h5fffdfff0, 48'h6fffefff1, 48'h1fffafff5, 48'hfffffffafffc, 48'h200010004, 48'h40001fffe, 48'h6fffffff7, 48'h80001fff4, 48'ha0003fff7, 48'hfffefffafff4, 48'hffedffedffec, 48'hffe7ffe9ffeb, 48'hfff5fff7fff8, 48'h600080009, 48'hd000e000f, 48'h600060005, 48'hfffefffcfff7, 48'hfffffffbfff3, 48'h5fffefff3, 48'h9fffffff2, 48'h8fffefff2, 48'hfffffff9fff2, 48'hfffafff8fff6, 48'hfffcfffeffff, 48'hffff00010003, 48'hffffffff0002, 48'hfffafffafff9, 48'hfffffffefffb, 48'hfff6fff5fff8, 48'hffeaffebffe9, 48'hfffaffed, 48'h6fffdffee, 48'h4fffcffed, 48'h6fffdffed, 48'h9fffdfff0, 48'hfff8fff4, 48'hfffafffaffff, 48'h100020004, 48'h60002ffff, 48'h50000fff8, 48'hfffcfff8fff2, 48'hffeeffecffed, 48'hfff1fff3fff5, 48'h200030004, 48'ha000b000b, 48'h800080006, 48'h1fffffffa, 48'hfffffffafff2, 48'h5fffdfff0, 48'h8fffffff1, 48'h9ffffffef, 48'h8fffdffed, 48'h9fffeffed, 48'h8fffdfff0, 48'hfffafff2, 48'hfffdfffbfff9, 48'h2, 48'h200030004, 48'hfffdfffdfffe, 48'hfff8fff7fff5, 48'hfff9fff8fff5, 48'hfff6fff3ffeb, 48'hfffffff7ffe8, 48'h5fffbffeb, 48'h4fffaffe9, 48'h6fffaffe9, 48'h9fffcffeb, 48'h5fffcffee, 48'hfffafff7fff3, 48'hfffdfffcfffb, 48'h700040002, 48'hfffffffefffa, 48'hfff4fff4fff4, 48'hfffbfffafffd, 48'hfffffffffffe, 48'hfffffffd, 48'hfffdfff9, 48'hfffafff1, 48'h4fffbffee, 48'h8fffeffee, 48'h8fffeffee, 48'h8fffeffee, 48'h8fffdffed, 48'h8fffdffec, 48'h8fffdffec, 48'h8fffcffed, 48'h6fffbffed, 48'hfffffff8ffef, 48'hfffffffdfffa, 48'hfffe0000ffff, 48'hfff8fffcfff8, 48'hfffafff8fff8, 48'hfffcfff6ffed, 48'h2fff8ffe9, 48'h2fff6ffe6, 48'h5fff9ffe7, 48'h4fff8ffe6, 48'h5fff8ffe6, 48'h9fffaffe7, 48'h6fffcffe6, 48'h1fffaffeb, 48'hfffdfff7fff2, 48'hfffdfffafff9, 48'hfff5fff8fff8, 48'hfff3fff7fffa, 48'hffefffeffff2, 48'hfff4fff0ffeb, 48'hfffffff7ffec, 48'h4fffaffed, 48'h8fffcffec, 48'h9fffcffea, 48'h8fffcffea, 48'h7fffcffeb, 48'h7fffcffea, 48'h8fffbffe9, 48'h8fffbffe8, 48'h6fffaffe9, 48'h8fffaffe9, 48'hafffbffe6, 48'h6fff9ffe8, 48'hfffbfff5ffed, 48'hfff5fff7fff8, 48'hfff7fffcffff, 48'hfff8fff8fffb, 48'hfffcfff7ffec, 48'h4fff8ffe3, 48'h5fff8ffe5, 48'h4fff7ffe4, 48'h4fff6ffe2, 48'h5fff7ffe2, 48'h8fff9ffe5, 48'h6fffbffe1, 48'h6fffbffe4, 48'hfffcfff4ffeb, 48'hffebffe9ffe9, 48'hffe6ffe9ffe9, 48'hffe9ffebffee, 48'hfff2fff2fff4, 48'hfffbfff7fff0, 48'h7fffaffea, 48'hbfffcffe8, 48'hafffbffe6, 48'h6fffaffe7, 48'h5fff9ffe8, 48'h6fffaffe8, 48'h7fffaffe7, 48'h8fffaffe6, 48'h8fffaffe5, 48'h6fff9ffe6, 48'h8fff9ffe5, 48'hafff9ffe2, 48'h8fff9ffe3, 48'h1fff7ffe7, 48'hfff3ffefffed, 48'hfff1fff1fffc, 48'hfff3fff7fffa, 48'hfff8fff7fff2, 48'hfffefff6ffe4, 48'h3fff7ffe1, 48'h3fff5ffe1, 48'h3fff5ffe0, 48'h5fff6ffe0, 48'h5fff7ffe3, 48'h5fff8ffe1, 48'h8fff9ffe1, 48'hfffbfff2ffe5, 48'hffe1ffe1ffe2, 48'hffe0ffe2ffe2, 48'hffeeffedffeb, 48'hfffbfff9fffa, 48'hfffefffcfff8, 48'h1fff8ffeb, 48'h6fff8ffe6, 48'h9fff9ffe3, 48'h8fff9ffe3, 48'h5fff8ffe4, 48'h5fff8ffe4, 48'h6fff8ffe3, 48'h6fff8ffe3, 48'h7fff8ffe2, 48'h6fff8ffe2, 48'h6fff8ffe2, 48'h6fff7ffe1, 48'h6fff7ffe1, 48'h5fff7ffe1, 48'hfffffff3ffe6, 48'hfff3ffeeffee, 48'hffeeffeffff6, 48'hfff3fff4fff8, 48'hfffbfff5ffee, 48'hfffffff4ffdf, 48'h1fff4ffde, 48'h1fff4ffdd, 48'h3fff5ffdd, 48'h3fff5ffe1, 48'h4fff6ffe0, 48'h8fff7ffde, 48'hfff8fff0ffe3, 48'hffe0ffe1ffe3, 48'hffe7ffe7ffe4, 48'hfff7fff1ffe8, 48'hfffafff3ffec, 48'hfffdfff9fff4, 48'hfffbfff4, 48'h1fff6ffe7, 48'h7fff7ffe1, 48'h9fff8ffdf, 48'h7fff7ffe0, 48'h5fff7ffe1, 48'h5fff6ffe0, 48'h6fff6ffe0, 48'h6fff6ffe0, 48'h6fff6ffdf, 48'h5fff6ffdf, 48'h4fff5ffe0, 48'h4fff5ffdf, 48'h6fff5ffdd, 48'h6fff5ffdd, 48'hfffdfff4ffe0, 48'hfff0ffecffed, 48'hfff1ffeffff8, 48'hfffafff7fffa, 48'hfffefff4ffe4, 48'hfffffff2ffdd, 48'h1fff3ffdc, 48'h3fff4ffdb, 48'h3fff4ffdf, 48'h4fff5ffdd, 48'h7fff6ffdb, 48'hfff4ffedffe3, 48'hffdfffe1ffe3, 48'hffedffe9ffe2, 48'h2fff4ffe2, 48'h3fff4ffe0, 48'hfffffff4ffe5, 48'hfff7ffec, 48'h2fff5ffe4, 48'h6fff5ffde, 48'h6fff6ffdd, 48'h5fff5ffde, 48'h6fff5ffde, 48'h6fff5ffde, 48'h5fff5ffdd, 48'h5fff5ffdd, 48'h5fff4ffdd, 48'h5fff4ffdd, 48'h5fff4ffdd, 48'h5fff4ffdd, 48'h5fff4ffdd, 48'h5fff4ffdc, 48'h2fff5ffda, 48'hfffafff1ffe1, 48'hfff3ffecffed, 48'hfff8fff4fff3, 48'hfffefff4ffe7, 48'hfffefff1ffdd, 48'h2fff2ffda, 48'h4fff2ffda, 48'h3fff3ffdd, 48'h3fff3ffdb, 48'h5fff4ffda, 48'hfff4ffecffe0, 48'hffe6ffe4ffe0, 48'hfff4ffedffe1, 48'h4fff4ffdd, 48'h6fff5ffdc, 48'h1fff3ffdf, 48'hfff3ffe1, 48'h4fff4ffde, 48'h6fff4ffdc, 48'h4fff4ffdc, 48'h3fff4ffdd, 48'h5fff4ffdc, 48'h5fff4ffdc, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h4fff3ffdc, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h6fff2ffdc, 48'h5fff3ffd8, 48'h2fff2ffdb, 48'hfffdffefffe1, 48'hfffcfff1ffdf, 48'hfffefff1ffdd, 48'hfffffff1ffda, 48'h1fff1ffd8, 48'h2fff1ffd8, 48'h3fff2ffdb, 48'h4fff2ffda, 48'h5fff3ffda, 48'hfff9ffedffdd, 48'hfff2ffebffde, 48'hfffdfff2ffdf, 48'h5fff4ffda, 48'h6fff4ffd8, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h6fff3ffda, 48'h6fff4ffda, 48'h4fff3ffdb, 48'h3fff3ffdc, 48'h4fff3ffdb, 48'h4fff3ffdb, 48'h4fff2ffda, 48'h4fff2ffda, 48'h4fff2ffda, 48'h4fff3ffda, 48'h4fff2ffda, 48'h4fff2ffda, 48'h4fff2ffda, 48'h4fff1ffda, 48'h5fff2ffd7, 48'h4fff2ffd7, 48'h4fff1ffda, 48'h4fff1ffd7, 48'h2fff1ffd8, 48'hfff0ffd7, 48'hfff0ffd6, 48'hfff0ffd7, 48'h3fff1ffda, 48'h4fff1ffda, 48'h4fff1ffda, 48'hfff1ffdc, 48'hfffdfff1ffdd, 48'h1fff2ffdb, 48'h5fff3ffd8, 48'h6fff3ffd8, 48'h5fff3ffd8, 48'h5fff3ffd8, 48'h6fff3ffd8, 48'h5fff3ffd8, 48'h4fff2ffd9, 48'h3fff2ffda, 48'h4fff2ffd9, 48'h4fff2ffd9, 48'h4fff2ffd9, 48'h4fff2ffd9, 48'h4fff2ffd9, 48'h3fff2ffd8, 48'h3fff1ffd8, 48'h3fff1ffd8, 48'h3fff1ffd8, 48'h2fff1ffd7, 48'h1fff1ffd6, 48'h2fff1ffd8, 48'h3ffefffd9, 48'h3ffeeffd9, 48'h2ffefffd6, 48'hffefffd5, 48'hffffffeeffd5, 48'hffffffeeffd6, 48'h3fff0ffd7, 48'h4ffefffd8, 48'h2ffefffda, 48'h2fff1ffd9, 48'h2fff1ffd9, 48'h2fff1ffd9, 48'h4fff1ffd8, 48'h4fff2ffd8, 48'h4fff2ffd8, 48'h4fff2ffd7, 48'h4fff2ffd7, 48'h4fff1ffd8, 48'h4fff1ffd8, 48'h4fff1ffd8, 48'h3fff1ffd8, 48'h3fff1ffd8, 48'h3fff1ffd7, 48'h3fff1ffd7, 48'h3fff1ffd7, 48'h2fff0ffd7, 48'h2fff0ffd7, 48'h2fff0ffd7, 48'h2fff0ffd7, 48'h1fff0ffd6, 48'hffefffd7, 48'hffefffd7, 48'hffeeffd7, 48'hffedffd7, 48'hffedffd6, 48'hffffffedffd5, 48'hfffdffecffd5, 48'hffedffd5};

   reg         clock;
   reg 	       reset;
   reg 	       vld_in;
   wire        vld_out;
   wire [63:0][15:0] bits_out;

   reg [9:0]   img_cntr;
   reg [9:0]   img_cntr_out;
   wire        bits_out_correct;
   wire [47:0] curr_pixel;
   assign curr_pixel = airplane4_image[img_cntr];
   wire [2:0][15:0] in;
   assign in[0] = curr_pixel[15:0];
   assign in[1] = curr_pixel[31:16];
   assign in[2] = curr_pixel[47:32];
   assign bits_out_correct = ( bits_out == airplane4_conv1[img_cntr_out] );
   
conv_windower lyr1_conv (
.clock(clock),
.reset(reset),
.vld_in(vld_in),
.in(in),
.vld_out(vld_out),
.out( bits_out )
);

always #2 clock = ~clock;

always @(posedge clock)
  begin
     if ( vld_in )
       begin
	  img_cntr <= img_cntr + 1'h1;
       end
     if ( vld_out )
       begin
	  img_cntr_out <= img_cntr_out + 1'h1;
	  if ( bits_out_correct )
	    begin
	       $display("ASSERTION PASSED: %h == %h", bits_out, airplane4_conv1[img_cntr_out]);
	    end else begin
	       $display("ASSERTION FAILED: %h == %h", bits_out, airplane4_conv1[img_cntr_out]);
	    end
       end
  end
initial begin
   clock = 0;
   reset = 1;
   vld_in = 0;
   img_cntr = 0;
   img_cntr_out = 0;
   #32
   reset = 0;
   #32
   vld_in = 1;
   #4096
   vld_in = 0;
   #100
   vld_in = 1;
   #4096
   vld_in = 0;
   #100
   $finish;   
end

endmodule

